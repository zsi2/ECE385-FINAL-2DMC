module main_menu

(

	input [9:0] DrawX,DrawY,
	
	output [23:0] main_rgb
	
);

parameter bit [1:0] mc_rom [20399:0]='{


00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
01,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
10,
10,
10,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
01,
01,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
01,
01,
01,
01,
10,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00

};

parameter bit [1:0] button_rom [15999:0]='{

00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
01,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
10,
10,
10,
10,
10,
10,
10,
10,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
01,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
11,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00,
00



};

int rely,relx,rely1;

assign rely=DrawY-59;
assign relx=DrawX-119;
assign rely1=DrawY-211;
always_comb
begin

	if((DrawX>119)&&(DrawX<519)&&(DrawY>60)&&(DrawY<111)) //Minecraft
	begin
		if(mc_rom[rely*400+relx]==2'b00)
			main_rgb=24'hd2e6ff;
		else if (mc_rom[rely*400+relx]==2'b01)
			main_rgb=24'h000000;
		else
			main_rgb=24'h777777;
		
	end
	
	else if((DrawX>119)&&(DrawX<519)&&(DrawY>211)&&(DrawY<251))
	begin
		if(button_rom[rely1*400+relx]==2'b00)
			main_rgb=24'hd2e6ff;
		else if (button_rom[rely*400+relx]==2'b01)
			main_rgb=24'h000000;
		else
			main_rgb=24'h777777;
		
	end
	else
		main_rgb=24'hd2e6ff;
end

endmodule