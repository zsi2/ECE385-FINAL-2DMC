// vga_driver_with_framebuffer_soc.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module vga_driver_with_framebuffer_soc (
		input  wire        clk_clk,            //   clk.clk
		output wire        epcs_dclk,          //  epcs.dclk
		output wire        epcs_sce,           //      .sce
		output wire        epcs_sdo,           //      .sdo
		input  wire        epcs_data0,         //      .data0
		input  wire        reset_reset_n,      // reset.reset_n
		output wire [12:0] sdram_addr,         // sdram.addr
		output wire [1:0]  sdram_ba,           //      .ba
		output wire        sdram_cas_n,        //      .cas_n
		output wire        sdram_cke,          //      .cke
		output wire        sdram_cs_n,         //      .cs_n
		inout  wire [31:0] sdram_dq,           //      .dq
		output wire [3:0]  sdram_dqm,          //      .dqm
		output wire        sdram_ras_n,        //      .ras_n
		output wire        sdram_we_n,         //      .we_n
		output wire        vga_export_vga_clk, //   vga.export_vga_clk
		output wire        vga_export_vga_hs,  //      .export_vga_hs
		output wire        vga_export_vga_vs,  //      .export_vga_vs
		output wire        vga_export_vga_de,  //      .export_vga_de
		output wire [7:0]  vga_export_vga_r,   //      .export_vga_r
		output wire [7:0]  vga_export_vga_g,   //      .export_vga_g
		output wire [7:0]  vga_export_vga_b    //      .export_vga_b
	);

	wire         lcd_sgdma_out_valid;                                                    // lcd_sgdma:out_valid -> sgdma_ta:in_valid
	wire  [31:0] lcd_sgdma_out_data;                                                     // lcd_sgdma:out_data -> sgdma_ta:in_data
	wire         lcd_sgdma_out_ready;                                                    // sgdma_ta:in_ready -> lcd_sgdma:out_ready
	wire         lcd_sgdma_out_startofpacket;                                            // lcd_sgdma:out_startofpacket -> sgdma_ta:in_startofpacket
	wire         lcd_sgdma_out_endofpacket;                                              // lcd_sgdma:out_endofpacket -> sgdma_ta:in_endofpacket
	wire   [1:0] lcd_sgdma_out_empty;                                                    // lcd_sgdma:out_empty -> sgdma_ta:in_empty
	wire         sgdma_ta_out_valid;                                                     // sgdma_ta:out_valid -> fifo_0:avalonst_sink_valid
	wire  [31:0] sgdma_ta_out_data;                                                      // sgdma_ta:out_data -> fifo_0:avalonst_sink_data
	wire         sgdma_ta_out_ready;                                                     // fifo_0:avalonst_sink_ready -> sgdma_ta:out_ready
	wire         sgdma_ta_out_startofpacket;                                             // sgdma_ta:out_startofpacket -> fifo_0:avalonst_sink_startofpacket
	wire         sgdma_ta_out_endofpacket;                                               // sgdma_ta:out_endofpacket -> fifo_0:avalonst_sink_endofpacket
	wire   [1:0] sgdma_ta_out_empty;                                                     // sgdma_ta:out_empty -> fifo_0:avalonst_sink_empty
	wire         sdram_sgdma_pll_c0_clk;                                                 // sdram_sgdma_pll:c0 -> [epcs_flash_controller_0:clk, fifo_0:wrclock, irq_mapper:clk, jtag_uart_0:clk, lcd_sgdma:clk, mm_interconnect_0:sdram_sgdma_pll_c0_clk, nios2_gen2_0:clk, onchip_memory2_0:clk, rst_controller:clk, sdram:clk, sgdma_ta:clk, sysid_qsys_0:clock]
	wire         vga_pll_c0_clk;                                                         // vga_pll:c0 -> [avalon_st_adapter:in_clk_0_clk, avalon_st_adapter_001:in_clk_0_clk, fifo_0:rdclock, rst_controller_001:clk, vga:clk, vga_ta:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                      // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                   // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                   // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [27:0] nios2_gen2_0_data_master_address;                                       // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                    // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                          // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                                 // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                         // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                     // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] lcd_sgdma_descriptor_read_readdata;                                     // mm_interconnect_0:lcd_sgdma_descriptor_read_readdata -> lcd_sgdma:descriptor_read_readdata
	wire         lcd_sgdma_descriptor_read_waitrequest;                                  // mm_interconnect_0:lcd_sgdma_descriptor_read_waitrequest -> lcd_sgdma:descriptor_read_waitrequest
	wire  [31:0] lcd_sgdma_descriptor_read_address;                                      // lcd_sgdma:descriptor_read_address -> mm_interconnect_0:lcd_sgdma_descriptor_read_address
	wire         lcd_sgdma_descriptor_read_read;                                         // lcd_sgdma:descriptor_read_read -> mm_interconnect_0:lcd_sgdma_descriptor_read_read
	wire         lcd_sgdma_descriptor_read_readdatavalid;                                // mm_interconnect_0:lcd_sgdma_descriptor_read_readdatavalid -> lcd_sgdma:descriptor_read_readdatavalid
	wire         lcd_sgdma_descriptor_write_waitrequest;                                 // mm_interconnect_0:lcd_sgdma_descriptor_write_waitrequest -> lcd_sgdma:descriptor_write_waitrequest
	wire  [31:0] lcd_sgdma_descriptor_write_address;                                     // lcd_sgdma:descriptor_write_address -> mm_interconnect_0:lcd_sgdma_descriptor_write_address
	wire         lcd_sgdma_descriptor_write_write;                                       // lcd_sgdma:descriptor_write_write -> mm_interconnect_0:lcd_sgdma_descriptor_write_write
	wire  [31:0] lcd_sgdma_descriptor_write_writedata;                                   // lcd_sgdma:descriptor_write_writedata -> mm_interconnect_0:lcd_sgdma_descriptor_write_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                               // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                            // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [27:0] nios2_gen2_0_instruction_master_address;                                // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                   // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                          // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire  [31:0] lcd_sgdma_m_read_readdata;                                              // mm_interconnect_0:lcd_sgdma_m_read_readdata -> lcd_sgdma:m_read_readdata
	wire         lcd_sgdma_m_read_waitrequest;                                           // mm_interconnect_0:lcd_sgdma_m_read_waitrequest -> lcd_sgdma:m_read_waitrequest
	wire  [31:0] lcd_sgdma_m_read_address;                                               // lcd_sgdma:m_read_address -> mm_interconnect_0:lcd_sgdma_m_read_address
	wire         lcd_sgdma_m_read_read;                                                  // lcd_sgdma:m_read_read -> mm_interconnect_0:lcd_sgdma_m_read_read
	wire         lcd_sgdma_m_read_readdatavalid;                                         // mm_interconnect_0:lcd_sgdma_m_read_readdatavalid -> lcd_sgdma:m_read_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;               // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;            // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;              // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                  // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                   // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire         mm_interconnect_0_lcd_sgdma_csr_chipselect;                             // mm_interconnect_0:lcd_sgdma_csr_chipselect -> lcd_sgdma:csr_chipselect
	wire  [31:0] mm_interconnect_0_lcd_sgdma_csr_readdata;                               // lcd_sgdma:csr_readdata -> mm_interconnect_0:lcd_sgdma_csr_readdata
	wire   [3:0] mm_interconnect_0_lcd_sgdma_csr_address;                                // mm_interconnect_0:lcd_sgdma_csr_address -> lcd_sgdma:csr_address
	wire         mm_interconnect_0_lcd_sgdma_csr_read;                                   // mm_interconnect_0:lcd_sgdma_csr_read -> lcd_sgdma:csr_read
	wire         mm_interconnect_0_lcd_sgdma_csr_write;                                  // mm_interconnect_0:lcd_sgdma_csr_write -> lcd_sgdma:csr_write
	wire  [31:0] mm_interconnect_0_lcd_sgdma_csr_writedata;                              // mm_interconnect_0:lcd_sgdma_csr_writedata -> lcd_sgdma:csr_writedata
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;             // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;             // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                 // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;               // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect; // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_chipselect -> epcs_flash_controller_0:chipselect
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata;   // epcs_flash_controller_0:readdata -> mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address;    // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_address -> epcs_flash_controller_0:address
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read;       // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_read -> epcs_flash_controller_0:read_n
	wire         mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write;      // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_write -> epcs_flash_controller_0:write_n
	wire  [31:0] mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata;  // mm_interconnect_0:epcs_flash_controller_0_epcs_control_port_writedata -> epcs_flash_controller_0:writedata
	wire  [31:0] mm_interconnect_0_fifo_0_in_csr_readdata;                               // fifo_0:wrclk_control_slave_readdata -> mm_interconnect_0:fifo_0_in_csr_readdata
	wire   [2:0] mm_interconnect_0_fifo_0_in_csr_address;                                // mm_interconnect_0:fifo_0_in_csr_address -> fifo_0:wrclk_control_slave_address
	wire         mm_interconnect_0_fifo_0_in_csr_read;                                   // mm_interconnect_0:fifo_0_in_csr_read -> fifo_0:wrclk_control_slave_read
	wire         mm_interconnect_0_fifo_0_in_csr_write;                                  // mm_interconnect_0:fifo_0_in_csr_write -> fifo_0:wrclk_control_slave_write
	wire  [31:0] mm_interconnect_0_fifo_0_in_csr_writedata;                              // mm_interconnect_0:fifo_0_in_csr_writedata -> fifo_0:wrclk_control_slave_writedata
	wire  [31:0] mm_interconnect_0_sdram_sgdma_pll_pll_slave_readdata;                   // sdram_sgdma_pll:readdata -> mm_interconnect_0:sdram_sgdma_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_sgdma_pll_pll_slave_address;                    // mm_interconnect_0:sdram_sgdma_pll_pll_slave_address -> sdram_sgdma_pll:address
	wire         mm_interconnect_0_sdram_sgdma_pll_pll_slave_read;                       // mm_interconnect_0:sdram_sgdma_pll_pll_slave_read -> sdram_sgdma_pll:read
	wire         mm_interconnect_0_sdram_sgdma_pll_pll_slave_write;                      // mm_interconnect_0:sdram_sgdma_pll_pll_slave_write -> sdram_sgdma_pll:write
	wire  [31:0] mm_interconnect_0_sdram_sgdma_pll_pll_slave_writedata;                  // mm_interconnect_0:sdram_sgdma_pll_pll_slave_writedata -> sdram_sgdma_pll:writedata
	wire  [31:0] mm_interconnect_0_vga_pll_pll_slave_readdata;                           // vga_pll:readdata -> mm_interconnect_0:vga_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_vga_pll_pll_slave_address;                            // mm_interconnect_0:vga_pll_pll_slave_address -> vga_pll:address
	wire         mm_interconnect_0_vga_pll_pll_slave_read;                               // mm_interconnect_0:vga_pll_pll_slave_read -> vga_pll:read
	wire         mm_interconnect_0_vga_pll_pll_slave_write;                              // mm_interconnect_0:vga_pll_pll_slave_write -> vga_pll:write
	wire  [31:0] mm_interconnect_0_vga_pll_pll_slave_writedata;                          // mm_interconnect_0:vga_pll_pll_slave_writedata -> vga_pll:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                  // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                    // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                 // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                     // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                        // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                                  // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                               // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                       // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                                   // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                       // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                         // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                          // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                       // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                            // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                        // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                            // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         irq_mapper_receiver0_irq;                                               // lcd_sgdma:csr_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                               // fifo_0:wrclk_control_slave_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                               // epcs_flash_controller_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                               // jtag_uart_0:av_irq -> irq_mapper:receiver3_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                   // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         vga_ta_out_valid;                                                       // vga_ta:out_valid -> avalon_st_adapter:in_0_valid
	wire  [31:0] vga_ta_out_data;                                                        // vga_ta:out_data -> avalon_st_adapter:in_0_data
	wire         vga_ta_out_ready;                                                       // avalon_st_adapter:in_0_ready -> vga_ta:out_ready
	wire         vga_ta_out_startofpacket;                                               // vga_ta:out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         vga_ta_out_endofpacket;                                                 // vga_ta:out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire   [1:0] vga_ta_out_empty;                                                       // vga_ta:out_empty -> avalon_st_adapter:in_0_empty
	wire         avalon_st_adapter_out_0_valid;                                          // avalon_st_adapter:out_0_valid -> vga:valid_in
	wire  [31:0] avalon_st_adapter_out_0_data;                                           // avalon_st_adapter:out_0_data -> vga:data_in
	wire         avalon_st_adapter_out_0_ready;                                          // vga:ready_out -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                                  // avalon_st_adapter:out_0_startofpacket -> vga:sop_in
	wire         avalon_st_adapter_out_0_endofpacket;                                    // avalon_st_adapter:out_0_endofpacket -> vga:eop_in
	wire   [1:0] avalon_st_adapter_out_0_empty;                                          // avalon_st_adapter:out_0_empty -> vga:empty_in
	wire         fifo_0_out_valid;                                                       // fifo_0:avalonst_source_valid -> avalon_st_adapter_001:in_0_valid
	wire  [31:0] fifo_0_out_data;                                                        // fifo_0:avalonst_source_data -> avalon_st_adapter_001:in_0_data
	wire         fifo_0_out_ready;                                                       // avalon_st_adapter_001:in_0_ready -> fifo_0:avalonst_source_ready
	wire         fifo_0_out_startofpacket;                                               // fifo_0:avalonst_source_startofpacket -> avalon_st_adapter_001:in_0_startofpacket
	wire         fifo_0_out_endofpacket;                                                 // fifo_0:avalonst_source_endofpacket -> avalon_st_adapter_001:in_0_endofpacket
	wire   [1:0] fifo_0_out_empty;                                                       // fifo_0:avalonst_source_empty -> avalon_st_adapter_001:in_0_empty
	wire         avalon_st_adapter_001_out_0_valid;                                      // avalon_st_adapter_001:out_0_valid -> vga_ta:in_valid
	wire  [31:0] avalon_st_adapter_001_out_0_data;                                       // avalon_st_adapter_001:out_0_data -> vga_ta:in_data
	wire         avalon_st_adapter_001_out_0_ready;                                      // vga_ta:in_ready -> avalon_st_adapter_001:out_0_ready
	wire         avalon_st_adapter_001_out_0_startofpacket;                              // avalon_st_adapter_001:out_0_startofpacket -> vga_ta:in_startofpacket
	wire         avalon_st_adapter_001_out_0_endofpacket;                                // avalon_st_adapter_001:out_0_endofpacket -> vga_ta:in_endofpacket
	wire   [1:0] avalon_st_adapter_001_out_0_empty;                                      // avalon_st_adapter_001:out_0_empty -> vga_ta:in_empty
	wire         rst_controller_reset_out_reset;                                         // rst_controller:reset_out -> [epcs_flash_controller_0:reset_n, fifo_0:wrreset_n, irq_mapper:reset, jtag_uart_0:rst_n, lcd_sgdma:system_reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram:reset_n, sgdma_ta:reset_n, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                                     // rst_controller:reset_req -> [epcs_flash_controller_0:reset_req, nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                                 // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                     // rst_controller_001:reset_out -> [avalon_st_adapter:in_rst_0_reset, avalon_st_adapter_001:in_rst_0_reset, fifo_0:rdreset_n, vga:reset_n, vga_ta:reset_n]
	wire         rst_controller_002_reset_out_reset;                                     // rst_controller_002:reset_out -> [mm_interconnect_0:sdram_sgdma_pll_inclk_interface_reset_reset_bridge_in_reset_reset, sdram_sgdma_pll:reset, vga_pll:reset]

	vga_driver_with_framebuffer_soc_epcs_flash_controller_0 epcs_flash_controller_0 (
		.clk        (sdram_sgdma_pll_c0_clk),                                                 //               clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.reset_req  (rst_controller_reset_out_reset_req),                                     //                  .reset_req
		.address    (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address),    // epcs_control_port.address
		.chipselect (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect), //                  .chipselect
		.read_n     (~mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read),      //                  .read_n
		.readdata   (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata),   //                  .readdata
		.write_n    (~mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write),     //                  .write_n
		.writedata  (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata),  //                  .writedata
		.irq        (irq_mapper_receiver2_irq),                                               //               irq.irq
		.dclk       (epcs_dclk),                                                              //          external.export
		.sce        (epcs_sce),                                                               //                  .export
		.sdo        (epcs_sdo),                                                               //                  .export
		.data0      (epcs_data0)                                                              //                  .export
	);

	vga_driver_with_framebuffer_soc_fifo_0 fifo_0 (
		.wrclock                       (sdram_sgdma_pll_c0_clk),                    //    clk_in.clk
		.wrreset_n                     (~rst_controller_reset_out_reset),           //  reset_in.reset_n
		.rdclock                       (vga_pll_c0_clk),                            //   clk_out.clk
		.rdreset_n                     (~rst_controller_001_reset_out_reset),       // reset_out.reset_n
		.avalonst_sink_valid           (sgdma_ta_out_valid),                        //        in.valid
		.avalonst_sink_data            (sgdma_ta_out_data),                         //          .data
		.avalonst_sink_startofpacket   (sgdma_ta_out_startofpacket),                //          .startofpacket
		.avalonst_sink_endofpacket     (sgdma_ta_out_endofpacket),                  //          .endofpacket
		.avalonst_sink_empty           (sgdma_ta_out_empty),                        //          .empty
		.avalonst_sink_ready           (sgdma_ta_out_ready),                        //          .ready
		.avalonst_source_valid         (fifo_0_out_valid),                          //       out.valid
		.avalonst_source_data          (fifo_0_out_data),                           //          .data
		.avalonst_source_startofpacket (fifo_0_out_startofpacket),                  //          .startofpacket
		.avalonst_source_endofpacket   (fifo_0_out_endofpacket),                    //          .endofpacket
		.avalonst_source_empty         (fifo_0_out_empty),                          //          .empty
		.avalonst_source_ready         (fifo_0_out_ready),                          //          .ready
		.wrclk_control_slave_address   (mm_interconnect_0_fifo_0_in_csr_address),   //    in_csr.address
		.wrclk_control_slave_read      (mm_interconnect_0_fifo_0_in_csr_read),      //          .read
		.wrclk_control_slave_writedata (mm_interconnect_0_fifo_0_in_csr_writedata), //          .writedata
		.wrclk_control_slave_write     (mm_interconnect_0_fifo_0_in_csr_write),     //          .write
		.wrclk_control_slave_readdata  (mm_interconnect_0_fifo_0_in_csr_readdata),  //          .readdata
		.wrclk_control_slave_irq       (irq_mapper_receiver1_irq)                   //    in_irq.irq
	);

	vga_driver_with_framebuffer_soc_jtag_uart_0 jtag_uart_0 (
		.clk            (sdram_sgdma_pll_c0_clk),                                      //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver3_irq)                                     //               irq.irq
	);

	vga_driver_with_framebuffer_soc_lcd_sgdma lcd_sgdma (
		.clk                           (sdram_sgdma_pll_c0_clk),                     //              clk.clk
		.system_reset_n                (~rst_controller_reset_out_reset),            //            reset.reset_n
		.csr_chipselect                (mm_interconnect_0_lcd_sgdma_csr_chipselect), //              csr.chipselect
		.csr_address                   (mm_interconnect_0_lcd_sgdma_csr_address),    //                 .address
		.csr_read                      (mm_interconnect_0_lcd_sgdma_csr_read),       //                 .read
		.csr_write                     (mm_interconnect_0_lcd_sgdma_csr_write),      //                 .write
		.csr_writedata                 (mm_interconnect_0_lcd_sgdma_csr_writedata),  //                 .writedata
		.csr_readdata                  (mm_interconnect_0_lcd_sgdma_csr_readdata),   //                 .readdata
		.descriptor_read_readdata      (lcd_sgdma_descriptor_read_readdata),         //  descriptor_read.readdata
		.descriptor_read_readdatavalid (lcd_sgdma_descriptor_read_readdatavalid),    //                 .readdatavalid
		.descriptor_read_waitrequest   (lcd_sgdma_descriptor_read_waitrequest),      //                 .waitrequest
		.descriptor_read_address       (lcd_sgdma_descriptor_read_address),          //                 .address
		.descriptor_read_read          (lcd_sgdma_descriptor_read_read),             //                 .read
		.descriptor_write_waitrequest  (lcd_sgdma_descriptor_write_waitrequest),     // descriptor_write.waitrequest
		.descriptor_write_address      (lcd_sgdma_descriptor_write_address),         //                 .address
		.descriptor_write_write        (lcd_sgdma_descriptor_write_write),           //                 .write
		.descriptor_write_writedata    (lcd_sgdma_descriptor_write_writedata),       //                 .writedata
		.csr_irq                       (irq_mapper_receiver0_irq),                   //          csr_irq.irq
		.m_read_readdata               (lcd_sgdma_m_read_readdata),                  //           m_read.readdata
		.m_read_readdatavalid          (lcd_sgdma_m_read_readdatavalid),             //                 .readdatavalid
		.m_read_waitrequest            (lcd_sgdma_m_read_waitrequest),               //                 .waitrequest
		.m_read_address                (lcd_sgdma_m_read_address),                   //                 .address
		.m_read_read                   (lcd_sgdma_m_read_read),                      //                 .read
		.out_data                      (lcd_sgdma_out_data),                         //              out.data
		.out_valid                     (lcd_sgdma_out_valid),                        //                 .valid
		.out_ready                     (lcd_sgdma_out_ready),                        //                 .ready
		.out_endofpacket               (lcd_sgdma_out_endofpacket),                  //                 .endofpacket
		.out_startofpacket             (lcd_sgdma_out_startofpacket),                //                 .startofpacket
		.out_empty                     (lcd_sgdma_out_empty)                         //                 .empty
	);

	vga_driver_with_framebuffer_soc_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (sdram_sgdma_pll_c0_clk),                                     //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	vga_driver_with_framebuffer_soc_onchip_memory2_0 onchip_memory2_0 (
		.clk        (sdram_sgdma_pll_c0_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	vga_driver_with_framebuffer_soc_sdram sdram (
		.clk            (sdram_sgdma_pll_c0_clk),                   //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	vga_driver_with_framebuffer_soc_sdram_sgdma_pll sdram_sgdma_pll (
		.clk                (clk_clk),                                               //       inclk_interface.clk
		.reset              (rst_controller_002_reset_out_reset),                    // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_sgdma_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_sgdma_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_sgdma_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_sgdma_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_sgdma_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_sgdma_pll_c0_clk),                                //                    c0.clk
		.c1                 (),                                                      //                    c1.clk
		.scandone           (),                                                      //           (terminated)
		.scandataout        (),                                                      //           (terminated)
		.areset             (1'b0),                                                  //           (terminated)
		.locked             (),                                                      //           (terminated)
		.phasedone          (),                                                      //           (terminated)
		.phasecounterselect (4'b0000),                                               //           (terminated)
		.phaseupdown        (1'b0),                                                  //           (terminated)
		.phasestep          (1'b0),                                                  //           (terminated)
		.scanclk            (1'b0),                                                  //           (terminated)
		.scanclkena         (1'b0),                                                  //           (terminated)
		.scandata           (1'b0),                                                  //           (terminated)
		.configupdate       (1'b0)                                                   //           (terminated)
	);

	vga_driver_with_framebuffer_soc_sgdma_ta sgdma_ta (
		.clk               (sdram_sgdma_pll_c0_clk),          //   clk.clk
		.reset_n           (~rst_controller_reset_out_reset), // reset.reset_n
		.in_data           (lcd_sgdma_out_data),              //    in.data
		.in_valid          (lcd_sgdma_out_valid),             //      .valid
		.in_ready          (lcd_sgdma_out_ready),             //      .ready
		.in_startofpacket  (lcd_sgdma_out_startofpacket),     //      .startofpacket
		.in_endofpacket    (lcd_sgdma_out_endofpacket),       //      .endofpacket
		.in_empty          (lcd_sgdma_out_empty),             //      .empty
		.out_data          (sgdma_ta_out_data),               //   out.data
		.out_valid         (sgdma_ta_out_valid),              //      .valid
		.out_ready         (sgdma_ta_out_ready),              //      .ready
		.out_startofpacket (sgdma_ta_out_startofpacket),      //      .startofpacket
		.out_endofpacket   (sgdma_ta_out_endofpacket),        //      .endofpacket
		.out_empty         (sgdma_ta_out_empty)               //      .empty
	);

	vga_driver_with_framebuffer_soc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (sdram_sgdma_pll_c0_clk),                                //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	VGA_SINK #(
		.SYMBOLS_PER_BEAT (4),
		.BITS_PER_SYMBOL  (8),
		.READY_LATENCY    (0),
		.MAX_CHANNEL      (0),
		.H_DISP           (640),
		.H_FPORCH         (16),
		.H_SYNC           (96),
		.H_BPORCH         (48),
		.V_DISP           (480),
		.V_FPORCH         (10),
		.V_SYNC           (2),
		.V_BPORCH         (33)
	) vga (
		.ready_out (avalon_st_adapter_out_0_ready),         // avalon_streaming_sink.ready
		.valid_in  (avalon_st_adapter_out_0_valid),         //                      .valid
		.data_in   (avalon_st_adapter_out_0_data),          //                      .data
		.sop_in    (avalon_st_adapter_out_0_startofpacket), //                      .startofpacket
		.eop_in    (avalon_st_adapter_out_0_endofpacket),   //                      .endofpacket
		.empty_in  (avalon_st_adapter_out_0_empty),         //                      .empty
		.vga_clk   (vga_export_vga_clk),                    //           conduit_end.export_vga_clk
		.vga_hs    (vga_export_vga_hs),                     //                      .export_vga_hs
		.vga_vs    (vga_export_vga_vs),                     //                      .export_vga_vs
		.vga_de    (vga_export_vga_de),                     //                      .export_vga_de
		.vga_r     (vga_export_vga_r),                      //                      .export_vga_r
		.vga_g     (vga_export_vga_g),                      //                      .export_vga_g
		.vga_b     (vga_export_vga_b),                      //                      .export_vga_b
		.reset_n   (~rst_controller_001_reset_out_reset),   //                 reset.reset_n
		.clk       (vga_pll_c0_clk)                         //                 clock.clk
	);

	vga_driver_with_framebuffer_soc_vga_pll vga_pll (
		.clk                (clk_clk),                                       //       inclk_interface.clk
		.reset              (rst_controller_002_reset_out_reset),            // inclk_interface_reset.reset
		.read               (mm_interconnect_0_vga_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_vga_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_vga_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_vga_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_vga_pll_pll_slave_writedata), //                      .writedata
		.c0                 (vga_pll_c0_clk),                                //                    c0.clk
		.scandone           (),                                              //           (terminated)
		.scandataout        (),                                              //           (terminated)
		.areset             (1'b0),                                          //           (terminated)
		.locked             (),                                              //           (terminated)
		.phasedone          (),                                              //           (terminated)
		.phasecounterselect (4'b0000),                                       //           (terminated)
		.phaseupdown        (1'b0),                                          //           (terminated)
		.phasestep          (1'b0),                                          //           (terminated)
		.scanclk            (1'b0),                                          //           (terminated)
		.scanclkena         (1'b0),                                          //           (terminated)
		.scandata           (1'b0),                                          //           (terminated)
		.configupdate       (1'b0)                                           //           (terminated)
	);

	vga_driver_with_framebuffer_soc_sgdma_ta vga_ta (
		.clk               (vga_pll_c0_clk),                            //   clk.clk
		.reset_n           (~rst_controller_001_reset_out_reset),       // reset.reset_n
		.in_data           (avalon_st_adapter_001_out_0_data),          //    in.data
		.in_valid          (avalon_st_adapter_001_out_0_valid),         //      .valid
		.in_ready          (avalon_st_adapter_001_out_0_ready),         //      .ready
		.in_startofpacket  (avalon_st_adapter_001_out_0_startofpacket), //      .startofpacket
		.in_endofpacket    (avalon_st_adapter_001_out_0_endofpacket),   //      .endofpacket
		.in_empty          (avalon_st_adapter_001_out_0_empty),         //      .empty
		.out_data          (vga_ta_out_data),                           //   out.data
		.out_valid         (vga_ta_out_valid),                          //      .valid
		.out_ready         (vga_ta_out_ready),                          //      .ready
		.out_startofpacket (vga_ta_out_startofpacket),                  //      .startofpacket
		.out_endofpacket   (vga_ta_out_endofpacket),                    //      .endofpacket
		.out_empty         (vga_ta_out_empty)                           //      .empty
	);

	vga_driver_with_framebuffer_soc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                     (clk_clk),                                                                //                                                   clk_0_clk.clk
		.sdram_sgdma_pll_c0_clk                                            (sdram_sgdma_pll_c0_clk),                                                 //                                          sdram_sgdma_pll_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset                    (rst_controller_reset_out_reset),                                         //                    nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.sdram_sgdma_pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                                     // sdram_sgdma_pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.lcd_sgdma_descriptor_read_address                                 (lcd_sgdma_descriptor_read_address),                                      //                                   lcd_sgdma_descriptor_read.address
		.lcd_sgdma_descriptor_read_waitrequest                             (lcd_sgdma_descriptor_read_waitrequest),                                  //                                                            .waitrequest
		.lcd_sgdma_descriptor_read_read                                    (lcd_sgdma_descriptor_read_read),                                         //                                                            .read
		.lcd_sgdma_descriptor_read_readdata                                (lcd_sgdma_descriptor_read_readdata),                                     //                                                            .readdata
		.lcd_sgdma_descriptor_read_readdatavalid                           (lcd_sgdma_descriptor_read_readdatavalid),                                //                                                            .readdatavalid
		.lcd_sgdma_descriptor_write_address                                (lcd_sgdma_descriptor_write_address),                                     //                                  lcd_sgdma_descriptor_write.address
		.lcd_sgdma_descriptor_write_waitrequest                            (lcd_sgdma_descriptor_write_waitrequest),                                 //                                                            .waitrequest
		.lcd_sgdma_descriptor_write_write                                  (lcd_sgdma_descriptor_write_write),                                       //                                                            .write
		.lcd_sgdma_descriptor_write_writedata                              (lcd_sgdma_descriptor_write_writedata),                                   //                                                            .writedata
		.lcd_sgdma_m_read_address                                          (lcd_sgdma_m_read_address),                                               //                                            lcd_sgdma_m_read.address
		.lcd_sgdma_m_read_waitrequest                                      (lcd_sgdma_m_read_waitrequest),                                           //                                                            .waitrequest
		.lcd_sgdma_m_read_read                                             (lcd_sgdma_m_read_read),                                                  //                                                            .read
		.lcd_sgdma_m_read_readdata                                         (lcd_sgdma_m_read_readdata),                                              //                                                            .readdata
		.lcd_sgdma_m_read_readdatavalid                                    (lcd_sgdma_m_read_readdatavalid),                                         //                                                            .readdatavalid
		.nios2_gen2_0_data_master_address                                  (nios2_gen2_0_data_master_address),                                       //                                    nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                              (nios2_gen2_0_data_master_waitrequest),                                   //                                                            .waitrequest
		.nios2_gen2_0_data_master_byteenable                               (nios2_gen2_0_data_master_byteenable),                                    //                                                            .byteenable
		.nios2_gen2_0_data_master_read                                     (nios2_gen2_0_data_master_read),                                          //                                                            .read
		.nios2_gen2_0_data_master_readdata                                 (nios2_gen2_0_data_master_readdata),                                      //                                                            .readdata
		.nios2_gen2_0_data_master_readdatavalid                            (nios2_gen2_0_data_master_readdatavalid),                                 //                                                            .readdatavalid
		.nios2_gen2_0_data_master_write                                    (nios2_gen2_0_data_master_write),                                         //                                                            .write
		.nios2_gen2_0_data_master_writedata                                (nios2_gen2_0_data_master_writedata),                                     //                                                            .writedata
		.nios2_gen2_0_data_master_debugaccess                              (nios2_gen2_0_data_master_debugaccess),                                   //                                                            .debugaccess
		.nios2_gen2_0_instruction_master_address                           (nios2_gen2_0_instruction_master_address),                                //                             nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                            //                                                            .waitrequest
		.nios2_gen2_0_instruction_master_read                              (nios2_gen2_0_instruction_master_read),                                   //                                                            .read
		.nios2_gen2_0_instruction_master_readdata                          (nios2_gen2_0_instruction_master_readdata),                               //                                                            .readdata
		.nios2_gen2_0_instruction_master_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),                          //                                                            .readdatavalid
		.epcs_flash_controller_0_epcs_control_port_address                 (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_address),    //                   epcs_flash_controller_0_epcs_control_port.address
		.epcs_flash_controller_0_epcs_control_port_write                   (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_write),      //                                                            .write
		.epcs_flash_controller_0_epcs_control_port_read                    (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_read),       //                                                            .read
		.epcs_flash_controller_0_epcs_control_port_readdata                (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_readdata),   //                                                            .readdata
		.epcs_flash_controller_0_epcs_control_port_writedata               (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_writedata),  //                                                            .writedata
		.epcs_flash_controller_0_epcs_control_port_chipselect              (mm_interconnect_0_epcs_flash_controller_0_epcs_control_port_chipselect), //                                                            .chipselect
		.fifo_0_in_csr_address                                             (mm_interconnect_0_fifo_0_in_csr_address),                                //                                               fifo_0_in_csr.address
		.fifo_0_in_csr_write                                               (mm_interconnect_0_fifo_0_in_csr_write),                                  //                                                            .write
		.fifo_0_in_csr_read                                                (mm_interconnect_0_fifo_0_in_csr_read),                                   //                                                            .read
		.fifo_0_in_csr_readdata                                            (mm_interconnect_0_fifo_0_in_csr_readdata),                               //                                                            .readdata
		.fifo_0_in_csr_writedata                                           (mm_interconnect_0_fifo_0_in_csr_writedata),                              //                                                            .writedata
		.jtag_uart_0_avalon_jtag_slave_address                             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                //                               jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                  //                                                            .write
		.jtag_uart_0_avalon_jtag_slave_read                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                   //                                                            .read
		.jtag_uart_0_avalon_jtag_slave_readdata                            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),               //                                                            .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),              //                                                            .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),            //                                                            .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),             //                                                            .chipselect
		.lcd_sgdma_csr_address                                             (mm_interconnect_0_lcd_sgdma_csr_address),                                //                                               lcd_sgdma_csr.address
		.lcd_sgdma_csr_write                                               (mm_interconnect_0_lcd_sgdma_csr_write),                                  //                                                            .write
		.lcd_sgdma_csr_read                                                (mm_interconnect_0_lcd_sgdma_csr_read),                                   //                                                            .read
		.lcd_sgdma_csr_readdata                                            (mm_interconnect_0_lcd_sgdma_csr_readdata),                               //                                                            .readdata
		.lcd_sgdma_csr_writedata                                           (mm_interconnect_0_lcd_sgdma_csr_writedata),                              //                                                            .writedata
		.lcd_sgdma_csr_chipselect                                          (mm_interconnect_0_lcd_sgdma_csr_chipselect),                             //                                                            .chipselect
		.nios2_gen2_0_debug_mem_slave_address                              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                 //                                nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                   //                                                            .write
		.nios2_gen2_0_debug_mem_slave_read                                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                    //                                                            .read
		.nios2_gen2_0_debug_mem_slave_readdata                             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),                //                                                            .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),               //                                                            .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),              //                                                            .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),             //                                                            .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),             //                                                            .debugaccess
		.onchip_memory2_0_s1_address                                       (mm_interconnect_0_onchip_memory2_0_s1_address),                          //                                         onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                         (mm_interconnect_0_onchip_memory2_0_s1_write),                            //                                                            .write
		.onchip_memory2_0_s1_readdata                                      (mm_interconnect_0_onchip_memory2_0_s1_readdata),                         //                                                            .readdata
		.onchip_memory2_0_s1_writedata                                     (mm_interconnect_0_onchip_memory2_0_s1_writedata),                        //                                                            .writedata
		.onchip_memory2_0_s1_byteenable                                    (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                       //                                                            .byteenable
		.onchip_memory2_0_s1_chipselect                                    (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                       //                                                            .chipselect
		.onchip_memory2_0_s1_clken                                         (mm_interconnect_0_onchip_memory2_0_s1_clken),                            //                                                            .clken
		.sdram_s1_address                                                  (mm_interconnect_0_sdram_s1_address),                                     //                                                    sdram_s1.address
		.sdram_s1_write                                                    (mm_interconnect_0_sdram_s1_write),                                       //                                                            .write
		.sdram_s1_read                                                     (mm_interconnect_0_sdram_s1_read),                                        //                                                            .read
		.sdram_s1_readdata                                                 (mm_interconnect_0_sdram_s1_readdata),                                    //                                                            .readdata
		.sdram_s1_writedata                                                (mm_interconnect_0_sdram_s1_writedata),                                   //                                                            .writedata
		.sdram_s1_byteenable                                               (mm_interconnect_0_sdram_s1_byteenable),                                  //                                                            .byteenable
		.sdram_s1_readdatavalid                                            (mm_interconnect_0_sdram_s1_readdatavalid),                               //                                                            .readdatavalid
		.sdram_s1_waitrequest                                              (mm_interconnect_0_sdram_s1_waitrequest),                                 //                                                            .waitrequest
		.sdram_s1_chipselect                                               (mm_interconnect_0_sdram_s1_chipselect),                                  //                                                            .chipselect
		.sdram_sgdma_pll_pll_slave_address                                 (mm_interconnect_0_sdram_sgdma_pll_pll_slave_address),                    //                                   sdram_sgdma_pll_pll_slave.address
		.sdram_sgdma_pll_pll_slave_write                                   (mm_interconnect_0_sdram_sgdma_pll_pll_slave_write),                      //                                                            .write
		.sdram_sgdma_pll_pll_slave_read                                    (mm_interconnect_0_sdram_sgdma_pll_pll_slave_read),                       //                                                            .read
		.sdram_sgdma_pll_pll_slave_readdata                                (mm_interconnect_0_sdram_sgdma_pll_pll_slave_readdata),                   //                                                            .readdata
		.sdram_sgdma_pll_pll_slave_writedata                               (mm_interconnect_0_sdram_sgdma_pll_pll_slave_writedata),                  //                                                            .writedata
		.sysid_qsys_0_control_slave_address                                (mm_interconnect_0_sysid_qsys_0_control_slave_address),                   //                                  sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                               (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                  //                                                            .readdata
		.vga_pll_pll_slave_address                                         (mm_interconnect_0_vga_pll_pll_slave_address),                            //                                           vga_pll_pll_slave.address
		.vga_pll_pll_slave_write                                           (mm_interconnect_0_vga_pll_pll_slave_write),                              //                                                            .write
		.vga_pll_pll_slave_read                                            (mm_interconnect_0_vga_pll_pll_slave_read),                               //                                                            .read
		.vga_pll_pll_slave_readdata                                        (mm_interconnect_0_vga_pll_pll_slave_readdata),                           //                                                            .readdata
		.vga_pll_pll_slave_writedata                                       (mm_interconnect_0_vga_pll_pll_slave_writedata)                           //                                                            .writedata
	);

	vga_driver_with_framebuffer_soc_irq_mapper irq_mapper (
		.clk           (sdram_sgdma_pll_c0_clk),         //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	vga_driver_with_framebuffer_soc_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (vga_pll_c0_clk),                        // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),    // in_rst_0.reset
		.in_0_data           (vga_ta_out_data),                       //     in_0.data
		.in_0_valid          (vga_ta_out_valid),                      //         .valid
		.in_0_ready          (vga_ta_out_ready),                      //         .ready
		.in_0_startofpacket  (vga_ta_out_startofpacket),              //         .startofpacket
		.in_0_endofpacket    (vga_ta_out_endofpacket),                //         .endofpacket
		.in_0_empty          (vga_ta_out_empty),                      //         .empty
		.out_0_data          (avalon_st_adapter_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_out_0_empty)          //         .empty
	);

	vga_driver_with_framebuffer_soc_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (1),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter_001 (
		.in_clk_0_clk        (vga_pll_c0_clk),                            // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_001_reset_out_reset),        // in_rst_0.reset
		.in_0_data           (fifo_0_out_data),                           //     in_0.data
		.in_0_valid          (fifo_0_out_valid),                          //         .valid
		.in_0_ready          (fifo_0_out_ready),                          //         .ready
		.in_0_startofpacket  (fifo_0_out_startofpacket),                  //         .startofpacket
		.in_0_endofpacket    (fifo_0_out_endofpacket),                    //         .endofpacket
		.in_0_empty          (fifo_0_out_empty),                          //         .empty
		.out_0_data          (avalon_st_adapter_001_out_0_data),          //    out_0.data
		.out_0_valid         (avalon_st_adapter_001_out_0_valid),         //         .valid
		.out_0_ready         (avalon_st_adapter_001_out_0_ready),         //         .ready
		.out_0_startofpacket (avalon_st_adapter_001_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_001_out_0_endofpacket),   //         .endofpacket
		.out_0_empty         (avalon_st_adapter_001_out_0_empty)          //         .empty
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_sgdma_pll_c0_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (vga_pll_c0_clk),                         //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
