module artrom
(
	input logic [3:0] id,
	
	input logic [5:0] relx,rely,
	
	input logic [6:0] steve_relx,steve_rely,
	
	
	output logic [23:0] rgb,steve_rgb
	

	
);
	parameter bit [23:0] rom_bedrock [1599:0]='{
	
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757


		
};

parameter bit [23:0] rom_wood [1599:0]='{

24'h463926,
24'h463926,
24'h695433,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h685332,
24'h685332,
24'h685332,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6d5837,
24'h6d5837,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h463926,
24'h463926,
24'h695433,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h685332,
24'h685332,
24'h685332,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6d5837,
24'h6d5837,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h6f5a39,
24'h6f5a39,
24'h382b18,
24'h382b18,
24'h382b18,
24'h3f321f,
24'h3f321f,
24'h987849,
24'h987849,
24'h987849,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h665130,
24'h99794a,
24'h99794a,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h685332,
24'h685332,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h957546,
24'h957546,
24'h957546,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h6f5a39,
24'h6f5a39,
24'h382b18,
24'h382b18,
24'h382b18,
24'h3f321f,
24'h3f321f,
24'h987849,
24'h987849,
24'h987849,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h665130,
24'h99794a,
24'h99794a,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h685332,
24'h685332,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h957546,
24'h957546,
24'h957546,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h6f5a39,
24'h6f5a39,
24'h382b18,
24'h382b18,
24'h382b18,
24'h3f321f,
24'h3f321f,
24'h987849,
24'h987849,
24'h987849,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h665130,
24'h99794a,
24'h99794a,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h685332,
24'h685332,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h957546,
24'h957546,
24'h957546,
24'h3a2d1a,
24'h3a2d1a,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h644f2e,
24'h644f2e,
24'h413421,
24'h413421,
24'h413421,
24'h685332,
24'h685332,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3e311e,
24'h3e311e,
24'h675231,
24'h675231,
24'h675231,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3a2d1a,
24'h3a2d1a,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h644f2e,
24'h644f2e,
24'h413421,
24'h413421,
24'h413421,
24'h685332,
24'h685332,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3e311e,
24'h3e311e,
24'h675231,
24'h675231,
24'h675231,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h99794a,
24'h99794a,
24'h99794a,
24'h6d5837,
24'h6d5837,
24'h453825,
24'h453825,
24'h453825,
24'h634e2d,
24'h634e2d,
24'h403320,
24'h403320,
24'h403320,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h987849,
24'h3d301d,
24'h3d301d,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h423522,
24'h423522,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6d5837,
24'h6d5837,
24'h453825,
24'h453825,
24'h453825,
24'h634e2d,
24'h634e2d,
24'h403320,
24'h403320,
24'h403320,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h987849,
24'h3d301d,
24'h3d301d,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h423522,
24'h423522,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6d5837,
24'h6d5837,
24'h453825,
24'h453825,
24'h453825,
24'h634e2d,
24'h634e2d,
24'h403320,
24'h403320,
24'h403320,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h987849,
24'h3d301d,
24'h3d301d,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h423522,
24'h423522,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6a5534,
24'h6a5534,
24'h413421,
24'h413421,
24'h413421,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h675231,
24'h6e5938,
24'h6e5938,
24'h423522,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3c2f1c,
24'h3c2f1c,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6a5534,
24'h6a5534,
24'h413421,
24'h413421,
24'h413421,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h675231,
24'h6e5938,
24'h6e5938,
24'h423522,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3c2f1c,
24'h3c2f1c,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6c5736,
24'h6c5736,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h665130,
24'h665130,
24'h665130,
24'h9a7a4b,
24'h9a7a4b,
24'h685332,
24'h685332,
24'h685332,
24'h665130,
24'h665130,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6b5635,
24'h6b5635,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h695433,
24'h695433,
24'h8f6f40,
24'h8f6f40,
24'h8f6f40,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h675231,
24'h675231,
24'h675231,
24'h6c5736,
24'h6c5736,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h665130,
24'h665130,
24'h665130,
24'h9a7a4b,
24'h9a7a4b,
24'h685332,
24'h685332,
24'h685332,
24'h665130,
24'h665130,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6b5635,
24'h6b5635,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h695433,
24'h695433,
24'h8f6f40,
24'h8f6f40,
24'h8f6f40,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h675231,
24'h675231,
24'h675231,
24'h6c5736,
24'h6c5736,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h665130,
24'h665130,
24'h665130,
24'h9a7a4b,
24'h9a7a4b,
24'h685332,
24'h685332,
24'h685332,
24'h665130,
24'h665130,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6b5635,
24'h6b5635,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h695433,
24'h695433,
24'h8f6f40,
24'h8f6f40,
24'h8f6f40,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h675231,
24'h675231,
24'h675231,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h624d2c,
24'h624d2c,
24'h624d2c,
24'h685332,
24'h685332,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h917142,
24'h917142,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h7c623e,
24'h7c623e,
24'h59472c,
24'h59472c,
24'h59472c,
24'h372a17,
24'h372a17,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h624d2c,
24'h624d2c,
24'h624d2c,
24'h685332,
24'h685332,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h917142,
24'h917142,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h7c623e,
24'h7c623e,
24'h59472c,
24'h59472c,
24'h59472c,
24'h372a17,
24'h372a17,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3e311e,
24'h3e311e,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h413421,
24'h413421,
24'h413421,
24'h99794a,
24'h99794a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h4c3d26,
24'h665130,
24'h665130,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3e311e,
24'h3e311e,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h413421,
24'h413421,
24'h413421,
24'h99794a,
24'h99794a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h4c3d26,
24'h665130,
24'h665130,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3e311e,
24'h3e311e,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h413421,
24'h413421,
24'h413421,
24'h99794a,
24'h99794a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h4c3d26,
24'h665130,
24'h665130,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h695433,
24'h695433,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3f321f,
24'h3f321f,
24'h705b3a,
24'h705b3a,
24'h705b3a,
24'h947445,
24'h947445,
24'h413421,
24'h413421,
24'h413421,
24'h695433,
24'h695433,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h423522,
24'h423522,
24'h423522,
24'h937344,
24'h937344,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h6c5736,
24'h6c5736,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h3f321f,
24'h3f321f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3f321f,
24'h3f321f,
24'h705b3a,
24'h705b3a,
24'h705b3a,
24'h947445,
24'h947445,
24'h413421,
24'h413421,
24'h413421,
24'h695433,
24'h695433,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h423522,
24'h423522,
24'h423522,
24'h937344,
24'h937344,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h6c5736,
24'h6c5736,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h3f321f,
24'h3f321f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h463926,
24'h463926,
24'h675231,
24'h675231,
24'h675231,
24'h6d5837,
24'h6d5837,
24'h947445,
24'h947445,
24'h947445,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h392c19,
24'h392c19,
24'h392c19,
24'h957546,
24'h957546,
24'h423522,
24'h423522,
24'h423522,
24'h6b5635,
24'h6b5635,
24'h957546,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h463926,
24'h463926,
24'h675231,
24'h675231,
24'h675231,
24'h6d5837,
24'h6d5837,
24'h947445,
24'h947445,
24'h947445,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h392c19,
24'h392c19,
24'h392c19,
24'h957546,
24'h957546,
24'h423522,
24'h423522,
24'h423522,
24'h6b5635,
24'h6b5635,
24'h957546,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h463926,
24'h463926,
24'h675231,
24'h675231,
24'h675231,
24'h6d5837,
24'h6d5837,
24'h947445,
24'h947445,
24'h947445,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h392c19,
24'h392c19,
24'h392c19,
24'h957546,
24'h957546,
24'h423522,
24'h423522,
24'h423522,
24'h6b5635,
24'h6b5635,
24'h957546,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h453825,
24'h453825,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h675231,
24'h675231,
24'h967647,
24'h967647,
24'h967647,
24'h3a2d1a,
24'h3a2d1a,
24'h644f2e,
24'h644f2e,
24'h644f2e,
24'h3e311e,
24'h3e311e,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9f7f50,
24'h9f7f50,
24'h403320,
24'h403320,
24'h403320,
24'h6a5534,
24'h6a5534,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h433623,
24'h433623,
24'h957546,
24'h957546,
24'h957546,
24'h453825,
24'h453825,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h675231,
24'h675231,
24'h967647,
24'h967647,
24'h967647,
24'h3a2d1a,
24'h3a2d1a,
24'h644f2e,
24'h644f2e,
24'h644f2e,
24'h3e311e,
24'h3e311e,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9f7f50,
24'h9f7f50,
24'h403320,
24'h403320,
24'h403320,
24'h6a5534,
24'h6a5534,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h433623,
24'h433623,
24'h957546,
24'h957546,
24'h957546,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h675231,
24'h675231,
24'h675231,
24'h6f5a39,
24'h6f5a39,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h423522,
24'h423522,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9d7d4e,
24'h9d7d4e,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h675231,
24'h675231,
24'h675231,
24'h6f5a39,
24'h6f5a39,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h423522,
24'h423522,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9d7d4e,
24'h9d7d4e,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h675231,
24'h675231,
24'h675231,
24'h6f5a39,
24'h6f5a39,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h423522,
24'h423522,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9d7d4e,
24'h9d7d4e,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3b2e1b,
24'h3b2e1b,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h392c19,
24'h392c19,
24'h665130,
24'h665130,
24'h665130,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h6a5534,
24'h6a5534,
24'h624d2c,
24'h624d2c,
24'h624d2c,
24'h403320,
24'h403320,
24'h987849,
24'h987849,
24'h987849,
24'h3b2e1b,
24'h3b2e1b,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h392c19,
24'h392c19,
24'h665130,
24'h665130,
24'h665130,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h6a5534,
24'h6a5534,
24'h624d2c,
24'h624d2c,
24'h624d2c,
24'h403320,
24'h403320,
24'h987849,
24'h987849,
24'h987849,
24'h413421,
24'h413421,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6d5837,
24'h6d5837,
24'h634e2d,
24'h634e2d,
24'h634e2d,
24'h675231,
24'h675231,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6a5534,
24'h6a5534,
24'h947445,
24'h947445,
24'h947445,
24'h9c7c4d,
24'h9c7c4d,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h413421,
24'h413421,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6d5837,
24'h6d5837,
24'h634e2d,
24'h634e2d,
24'h634e2d,
24'h675231,
24'h675231,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6a5534,
24'h6a5534,
24'h947445,
24'h947445,
24'h947445,
24'h9c7c4d,
24'h9c7c4d,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h413421,
24'h413421,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6d5837,
24'h6d5837,
24'h634e2d,
24'h634e2d,
24'h634e2d,
24'h675231,
24'h675231,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6a5534,
24'h6a5534,
24'h947445,
24'h947445,
24'h947445,
24'h9c7c4d,
24'h9c7c4d,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h675231,
24'h675231,
24'h675231,
24'h977748,
24'h977748,
24'h403320,
24'h403320,
24'h403320,
24'h6b5635,
24'h6b5635,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h927243,
24'h927243,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3b2e1b,
24'h3b2e1b,
24'h3b2e1b,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3d301d,
24'h3d301d,
24'h675231,
24'h675231,
24'h675231,
24'h3a2d1a,
24'h3a2d1a,
24'h675231,
24'h675231,
24'h675231,
24'h977748,
24'h977748,
24'h403320,
24'h403320,
24'h403320,
24'h6b5635,
24'h6b5635,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h927243,
24'h927243,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3b2e1b,
24'h3b2e1b,
24'h3b2e1b,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3d301d,
24'h3d301d,
24'h675231,
24'h675231,
24'h675231,
24'h5e4b2f,
24'h5e4b2f,
24'h685332,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h644f2e,
24'h644f2e,
24'h695433,
24'h695433,
24'h695433,
24'h685332,
24'h685332,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h372a17,
24'h372a17,
24'h372a17,
24'h675231,
24'h675231,
24'h695433,
24'h695433,
24'h695433,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h5e4b2f,
24'h5e4b2f,
24'h685332,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h644f2e,
24'h644f2e,
24'h695433,
24'h695433,
24'h695433,
24'h685332,
24'h685332,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h372a17,
24'h372a17,
24'h372a17,
24'h675231,
24'h675231,
24'h695433,
24'h695433,
24'h695433,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h5e4b2f,
24'h5e4b2f,
24'h685332,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h644f2e,
24'h644f2e,
24'h695433,
24'h695433,
24'h695433,
24'h685332,
24'h685332,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h372a17,
24'h372a17,
24'h372a17,
24'h675231,
24'h675231,
24'h695433,
24'h695433,
24'h695433,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e




};

parameter bit [23:0] rom_stone [1599:0]='{

24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h808080,
24'h808080,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h808080,
24'h808080,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h808080,
24'h808080,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f





};

parameter bit [23:0] rom_dirt [1599:0]='{


24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a




};

parameter bit [23:0] rom_steve [3199:0] ='{

24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h1b1004,
24'h1b1004,
24'h1b1004,
24'h170d01,
24'h170d01,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h100800,
24'h100800,
24'h0d0600,
24'h0d0600,
24'h0d0600,
24'h100800,
24'h100800,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h1b1004,
24'h1b1004,
24'h1b1004,
24'h170d01,
24'h170d01,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h100800,
24'h100800,
24'h0d0600,
24'h0d0600,
24'h0d0600,
24'h100800,
24'h100800,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h1b1004,
24'h1b1004,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h1b1004,
24'h1b1004,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h1b1004,
24'h1b1004,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h956f5a,
24'h956f5a,
24'h936551,
24'h936551,
24'h936551,
24'h946b57,
24'h946b57,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h211508,
24'h211508,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h956f5a,
24'h956f5a,
24'h936551,
24'h936551,
24'h936551,
24'h946b57,
24'h946b57,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h211508,
24'h211508,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h956f5a,
24'h956f5a,
24'h936551,
24'h936551,
24'h936551,
24'h946b57,
24'h946b57,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h211508,
24'h211508,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h915c48,
24'h915c48,
24'h915c48,
24'h946752,
24'h946752,
24'h915c48,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h936551,
24'h936551,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h915c48,
24'h915c48,
24'h915c48,
24'h946752,
24'h946752,
24'h915c48,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h936551,
24'h936551,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h946752,
24'h946752,
24'h946752,
24'hffffff,
24'hffffff,
24'h312877,
24'h312877,
24'h312877,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h312877,
24'h312877,
24'hffffff,
24'hffffff,
24'hffffff,
24'h915c48,
24'h915c48,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h946752,
24'h946752,
24'h946752,
24'hffffff,
24'hffffff,
24'h312877,
24'h312877,
24'h312877,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h312877,
24'h312877,
24'hffffff,
24'hffffff,
24'hffffff,
24'h915c48,
24'h915c48,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h7b4435,
24'h7b4435,
24'h7b4435,
24'h8b5441,
24'h8b5441,
24'h936551,
24'h936551,
24'h936551,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h936551,
24'h936551,
24'h8d5441,
24'h8d5441,
24'h8d5441,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h7b4435,
24'h7b4435,
24'h7b4435,
24'h8b5441,
24'h8b5441,
24'h936551,
24'h936551,
24'h936551,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h936551,
24'h936551,
24'h8d5441,
24'h8d5441,
24'h8d5441,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h7b4435,
24'h7b4435,
24'h7b4435,
24'h8b5441,
24'h8b5441,
24'h936551,
24'h936551,
24'h936551,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h936551,
24'h936551,
24'h8d5441,
24'h8d5441,
24'h8d5441,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h7b4435,
24'h7b4435,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h713b2d,
24'h713b2d,
24'h713b2d,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h7b4435,
24'h7b4435,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h713b2d,
24'h713b2d,
24'h713b2d,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h7b4435,
24'h7b4435,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h713b2d,
24'h713b2d,
24'h713b2d,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h764031,
24'h764031,
24'h764031,
24'h764031,
24'h764031,
24'h6a3a2d,
24'h6a3a2d,
24'h6a3a2d,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h60362c,
24'h60362c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h764031,
24'h764031,
24'h764031,
24'h764031,
24'h764031,
24'h6a3a2d,
24'h6a3a2d,
24'h6a3a2d,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h60362c,
24'h60362c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h905944,
24'h905944,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h905944,
24'h905944,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff



};

	
parameter bit [23:0] rom_diamond_ore[1599:0]
='{24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'hffffff,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h5decf5,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797
};
parameter bit [23:0] rom_furnace[1599:0]
='{24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757
};
parameter bit [23:0] rom_gold_ore[1599:0]
='{24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hffffff,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hffffff,
24'hffffff,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'hfcee4b,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797
};
parameter bit [23:0] rom_grass[1599:0]
='{24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a
};
parameter bit [23:0] rom_iron_ore[1599:0]
='{24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797
};
parameter bit [23:0] rom_leaves[1599:0]
='{24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813,
24'h00f265,
24'h00f265,
24'h00f265,
24'h3c9813,
24'h3c9813
};
parameter bit [23:0] rom_coal_ore[1599:0]
='{24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797
};
parameter bit [23:0] rom_crafting_table[1599:0]
='{24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h979797,
24'h979797,
24'h979797,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h433621,
24'h433621,
24'h433621,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h433621,
24'h000000,
24'h000000,
24'h000000
};
parameter bit [23:0] rom_water[1599:0]
='{24'h4c41f4,
24'h4c41f4,
24'h4633fe,
24'h4633fe,
24'h4633fe,
24'h363cff,
24'h363cff,
24'h4d32fc,
24'h4d32fc,
24'h4d32fc,
24'h4a2dff,
24'h4a2dff,
24'h3f32fd,
24'h3f32fd,
24'h3f32fd,
24'h4235ff,
24'h4235ff,
24'h4336ff,
24'h4336ff,
24'h4336ff,
24'h493cff,
24'h493cff,
24'h4235ff,
24'h4235ff,
24'h4235ff,
24'h4335ff,
24'h4335ff,
24'h4436ff,
24'h4436ff,
24'h4436ff,
24'h493bff,
24'h493bff,
24'h4c40f7,
24'h4c40f7,
24'h4c40f7,
24'h594bff,
24'h594bff,
24'h5241e6,
24'h5241e6,
24'h5241e6,
24'h4c41f4,
24'h4c41f4,
24'h4633fe,
24'h4633fe,
24'h4633fe,
24'h363cff,
24'h363cff,
24'h4d32fc,
24'h4d32fc,
24'h4d32fc,
24'h4a2dff,
24'h4a2dff,
24'h3f32fd,
24'h3f32fd,
24'h3f32fd,
24'h4235ff,
24'h4235ff,
24'h4336ff,
24'h4336ff,
24'h4336ff,
24'h493cff,
24'h493cff,
24'h4235ff,
24'h4235ff,
24'h4235ff,
24'h4335ff,
24'h4335ff,
24'h4436ff,
24'h4436ff,
24'h4436ff,
24'h493bff,
24'h493bff,
24'h4c40f7,
24'h4c40f7,
24'h4c40f7,
24'h594bff,
24'h594bff,
24'h5241e6,
24'h5241e6,
24'h5241e6,
24'h4c39ff,
24'h4c39ff,
24'h4f36ff,
24'h4f36ff,
24'h4f36ff,
24'h414afe,
24'h414afe,
24'h4841f2,
24'h4841f2,
24'h4841f2,
24'h4e4fff,
24'h4e4fff,
24'h4847fc,
24'h4847fc,
24'h4847fc,
24'h4c4bff,
24'h4c4bff,
24'h4745fd,
24'h4745fd,
24'h4745fd,
24'h4846fe,
24'h4846fe,
24'h4d4bff,
24'h4d4bff,
24'h4d4bff,
24'h4846ff,
24'h4846ff,
24'h3a38f2,
24'h3a38f2,
24'h3a38f2,
24'h4442fc,
24'h4442fc,
24'h473cff,
24'h473cff,
24'h473cff,
24'h3b2bff,
24'h3b2bff,
24'h4b36ff,
24'h4b36ff,
24'h4b36ff,
24'h4c39ff,
24'h4c39ff,
24'h4f36ff,
24'h4f36ff,
24'h4f36ff,
24'h414afe,
24'h414afe,
24'h4841f2,
24'h4841f2,
24'h4841f2,
24'h4e4fff,
24'h4e4fff,
24'h4847fc,
24'h4847fc,
24'h4847fc,
24'h4c4bff,
24'h4c4bff,
24'h4745fd,
24'h4745fd,
24'h4745fd,
24'h4846fe,
24'h4846fe,
24'h4d4bff,
24'h4d4bff,
24'h4d4bff,
24'h4846ff,
24'h4846ff,
24'h3a38f2,
24'h3a38f2,
24'h3a38f2,
24'h4442fc,
24'h4442fc,
24'h473cff,
24'h473cff,
24'h473cff,
24'h3b2bff,
24'h3b2bff,
24'h4b36ff,
24'h4b36ff,
24'h4b36ff,
24'h4c39ff,
24'h4c39ff,
24'h4f36ff,
24'h4f36ff,
24'h4f36ff,
24'h414afe,
24'h414afe,
24'h4841f2,
24'h4841f2,
24'h4841f2,
24'h4e4fff,
24'h4e4fff,
24'h4847fc,
24'h4847fc,
24'h4847fc,
24'h4c4bff,
24'h4c4bff,
24'h4745fd,
24'h4745fd,
24'h4745fd,
24'h4846fe,
24'h4846fe,
24'h4d4bff,
24'h4d4bff,
24'h4d4bff,
24'h4846ff,
24'h4846ff,
24'h3a38f2,
24'h3a38f2,
24'h3a38f2,
24'h4442fc,
24'h4442fc,
24'h473cff,
24'h473cff,
24'h473cff,
24'h3b2bff,
24'h3b2bff,
24'h4b36ff,
24'h4b36ff,
24'h4b36ff,
24'h3834fa,
24'h3834fa,
24'h3f35f7,
24'h3f35f7,
24'h3f35f7,
24'h3d3aff,
24'h3d3aff,
24'h4f36ff,
24'h4f36ff,
24'h4f36ff,
24'h4135f6,
24'h4135f6,
24'h4e44ff,
24'h4e44ff,
24'h4e44ff,
24'h4137f7,
24'h4137f7,
24'h4339f9,
24'h4339f9,
24'h4339f9,
24'h3e34f6,
24'h3e34f6,
24'h443afc,
24'h443afc,
24'h443afc,
24'h3f33f8,
24'h3f33f8,
24'h4d41ff,
24'h4d41ff,
24'h4d41ff,
24'h5044ff,
24'h5044ff,
24'h3c34fa,
24'h3c34fa,
24'h3c34fa,
24'h3f33f6,
24'h3f33f6,
24'h4a35fb,
24'h4a35fb,
24'h4a35fb,
24'h3834fa,
24'h3834fa,
24'h3f35f7,
24'h3f35f7,
24'h3f35f7,
24'h3d3aff,
24'h3d3aff,
24'h4f36ff,
24'h4f36ff,
24'h4f36ff,
24'h4135f6,
24'h4135f6,
24'h4e44ff,
24'h4e44ff,
24'h4e44ff,
24'h4137f7,
24'h4137f7,
24'h4339f9,
24'h4339f9,
24'h4339f9,
24'h3e34f6,
24'h3e34f6,
24'h443afc,
24'h443afc,
24'h443afc,
24'h3f33f8,
24'h3f33f8,
24'h4d41ff,
24'h4d41ff,
24'h4d41ff,
24'h5044ff,
24'h5044ff,
24'h3c34fa,
24'h3c34fa,
24'h3c34fa,
24'h3f33f6,
24'h3f33f6,
24'h4a35fb,
24'h4a35fb,
24'h4a35fb,
24'h4a39ff,
24'h4a39ff,
24'h4c41f6,
24'h4c41f6,
24'h4c41f6,
24'h5142ff,
24'h5142ff,
24'h4431fe,
24'h4431fe,
24'h4431fe,
24'h3c40f6,
24'h3c40f6,
24'h5347ff,
24'h5347ff,
24'h5347ff,
24'h4d41ff,
24'h4d41ff,
24'h5246ff,
24'h5246ff,
24'h5246ff,
24'h5244ff,
24'h5244ff,
24'h4739ff,
24'h4739ff,
24'h4739ff,
24'h4032fa,
24'h4032fa,
24'h4738ff,
24'h4738ff,
24'h4738ff,
24'h402ff9,
24'h402ff9,
24'h3d34f0,
24'h3d34f0,
24'h3d34f0,
24'h4a3ef9,
24'h4a3ef9,
24'h452ff5,
24'h452ff5,
24'h452ff5,
24'h4a39ff,
24'h4a39ff,
24'h4c41f6,
24'h4c41f6,
24'h4c41f6,
24'h5142ff,
24'h5142ff,
24'h4431fe,
24'h4431fe,
24'h4431fe,
24'h3c40f6,
24'h3c40f6,
24'h5347ff,
24'h5347ff,
24'h5347ff,
24'h4d41ff,
24'h4d41ff,
24'h5246ff,
24'h5246ff,
24'h5246ff,
24'h5244ff,
24'h5244ff,
24'h4739ff,
24'h4739ff,
24'h4739ff,
24'h4032fa,
24'h4032fa,
24'h4738ff,
24'h4738ff,
24'h4738ff,
24'h402ff9,
24'h402ff9,
24'h3d34f0,
24'h3d34f0,
24'h3d34f0,
24'h4a3ef9,
24'h4a3ef9,
24'h452ff5,
24'h452ff5,
24'h452ff5,
24'h4a39ff,
24'h4a39ff,
24'h4c41f6,
24'h4c41f6,
24'h4c41f6,
24'h5142ff,
24'h5142ff,
24'h4431fe,
24'h4431fe,
24'h4431fe,
24'h3c40f6,
24'h3c40f6,
24'h5347ff,
24'h5347ff,
24'h5347ff,
24'h4d41ff,
24'h4d41ff,
24'h5246ff,
24'h5246ff,
24'h5246ff,
24'h5244ff,
24'h5244ff,
24'h4739ff,
24'h4739ff,
24'h4739ff,
24'h4032fa,
24'h4032fa,
24'h4738ff,
24'h4738ff,
24'h4738ff,
24'h402ff9,
24'h402ff9,
24'h3d34f0,
24'h3d34f0,
24'h3d34f0,
24'h4a3ef9,
24'h4a3ef9,
24'h452ff5,
24'h452ff5,
24'h452ff5,
24'h4242ff,
24'h4242ff,
24'h3c4cff,
24'h3c4cff,
24'h3c4cff,
24'h504bff,
24'h504bff,
24'h4531ff,
24'h4531ff,
24'h4531ff,
24'h3a34ff,
24'h3a34ff,
24'h3a34f5,
24'h3a34f5,
24'h3a34f5,
24'h3e38f9,
24'h3e38f9,
24'h3d37f8,
24'h3d37f8,
24'h3d37f8,
24'h3f37fb,
24'h3f37fb,
24'h463eff,
24'h463eff,
24'h463eff,
24'h4139ff,
24'h4139ff,
24'h463bff,
24'h463bff,
24'h463bff,
24'h4136fe,
24'h4136fe,
24'h4335ff,
24'h4335ff,
24'h4335ff,
24'h4431ff,
24'h4431ff,
24'h4d33ff,
24'h4d33ff,
24'h4d33ff,
24'h4242ff,
24'h4242ff,
24'h3c4cff,
24'h3c4cff,
24'h3c4cff,
24'h504bff,
24'h504bff,
24'h4531ff,
24'h4531ff,
24'h4531ff,
24'h3a34ff,
24'h3a34ff,
24'h3a34f5,
24'h3a34f5,
24'h3a34f5,
24'h3e38f9,
24'h3e38f9,
24'h3d37f8,
24'h3d37f8,
24'h3d37f8,
24'h3f37fb,
24'h3f37fb,
24'h463eff,
24'h463eff,
24'h463eff,
24'h4139ff,
24'h4139ff,
24'h463bff,
24'h463bff,
24'h463bff,
24'h4136fe,
24'h4136fe,
24'h4335ff,
24'h4335ff,
24'h4335ff,
24'h4431ff,
24'h4431ff,
24'h4d33ff,
24'h4d33ff,
24'h4d33ff,
24'h4d48fc,
24'h4d48fc,
24'h4638fc,
24'h4638fc,
24'h4638fc,
24'h423bff,
24'h423bff,
24'h3d30ff,
24'h3d30ff,
24'h3d30ff,
24'h403af1,
24'h403af1,
24'h4634ff,
24'h4634ff,
24'h4634ff,
24'h4435ff,
24'h4435ff,
24'h473cff,
24'h473cff,
24'h473cff,
24'h4a3dff,
24'h4a3dff,
24'h4836ff,
24'h4836ff,
24'h4836ff,
24'h4632ff,
24'h4632ff,
24'h4232ff,
24'h4232ff,
24'h4232ff,
24'h3e30fe,
24'h3e30fe,
24'h4b47ff,
24'h4b47ff,
24'h4b47ff,
24'h4238fa,
24'h4238fa,
24'h4330fa,
24'h4330fa,
24'h4330fa,
24'h4d48fc,
24'h4d48fc,
24'h4638fc,
24'h4638fc,
24'h4638fc,
24'h423bff,
24'h423bff,
24'h3d30ff,
24'h3d30ff,
24'h3d30ff,
24'h403af1,
24'h403af1,
24'h4634ff,
24'h4634ff,
24'h4634ff,
24'h4435ff,
24'h4435ff,
24'h473cff,
24'h473cff,
24'h473cff,
24'h4a3dff,
24'h4a3dff,
24'h4836ff,
24'h4836ff,
24'h4836ff,
24'h4632ff,
24'h4632ff,
24'h4232ff,
24'h4232ff,
24'h4232ff,
24'h3e30fe,
24'h3e30fe,
24'h4b47ff,
24'h4b47ff,
24'h4b47ff,
24'h4238fa,
24'h4238fa,
24'h4330fa,
24'h4330fa,
24'h4330fa,
24'h4d48fc,
24'h4d48fc,
24'h4638fc,
24'h4638fc,
24'h4638fc,
24'h423bff,
24'h423bff,
24'h3d30ff,
24'h3d30ff,
24'h3d30ff,
24'h403af1,
24'h403af1,
24'h4634ff,
24'h4634ff,
24'h4634ff,
24'h4435ff,
24'h4435ff,
24'h473cff,
24'h473cff,
24'h473cff,
24'h4a3dff,
24'h4a3dff,
24'h4836ff,
24'h4836ff,
24'h4836ff,
24'h4632ff,
24'h4632ff,
24'h4232ff,
24'h4232ff,
24'h4232ff,
24'h3e30fe,
24'h3e30fe,
24'h4b47ff,
24'h4b47ff,
24'h4b47ff,
24'h4238fa,
24'h4238fa,
24'h4330fa,
24'h4330fa,
24'h4330fa,
24'h3c3cf1,
24'h3c3cf1,
24'h4c34fb,
24'h4c34fb,
24'h4c34fb,
24'h4131ff,
24'h4131ff,
24'h3e30ff,
24'h3e30ff,
24'h3e30ff,
24'h493dff,
24'h493dff,
24'h4636fa,
24'h4636fa,
24'h4636fa,
24'h453af9,
24'h453af9,
24'h483ffb,
24'h483ffb,
24'h483ffb,
24'h463bfa,
24'h463bfa,
24'h3e30f4,
24'h3e30f4,
24'h3e30f4,
24'h3f2ef5,
24'h3f2ef5,
24'h4337fa,
24'h4337fa,
24'h4337fa,
24'h463dfb,
24'h463dfb,
24'h4944ff,
24'h4944ff,
24'h4944ff,
24'h4d42ff,
24'h4d42ff,
24'h5946ff,
24'h5946ff,
24'h5946ff,
24'h3c3cf1,
24'h3c3cf1,
24'h4c34fb,
24'h4c34fb,
24'h4c34fb,
24'h4131ff,
24'h4131ff,
24'h3e30ff,
24'h3e30ff,
24'h3e30ff,
24'h493dff,
24'h493dff,
24'h4636fa,
24'h4636fa,
24'h4636fa,
24'h453af9,
24'h453af9,
24'h483ffb,
24'h483ffb,
24'h483ffb,
24'h463bfa,
24'h463bfa,
24'h3e30f4,
24'h3e30f4,
24'h3e30f4,
24'h3f2ef5,
24'h3f2ef5,
24'h4337fa,
24'h4337fa,
24'h4337fa,
24'h463dfb,
24'h463dfb,
24'h4944ff,
24'h4944ff,
24'h4944ff,
24'h4d42ff,
24'h4d42ff,
24'h5946ff,
24'h5946ff,
24'h5946ff,
24'h463aff,
24'h463aff,
24'h3b2ef6,
24'h3b2ef6,
24'h3b2ef6,
24'h4e4dff,
24'h4e4dff,
24'h4e47ff,
24'h4e47ff,
24'h4e47ff,
24'h4a3dee,
24'h4a3dee,
24'h4735ff,
24'h4735ff,
24'h4735ff,
24'h4235fd,
24'h4235fd,
24'h4237fc,
24'h4237fc,
24'h4237fc,
24'h4338fd,
24'h4338fd,
24'h4336ff,
24'h4336ff,
24'h4336ff,
24'h493aff,
24'h493aff,
24'h4e43ff,
24'h4e43ff,
24'h4e43ff,
24'h4d47ff,
24'h4d47ff,
24'h4540fd,
24'h4540fd,
24'h4540fd,
24'h4539fe,
24'h4539fe,
24'h422ffa,
24'h422ffa,
24'h422ffa,
24'h463aff,
24'h463aff,
24'h3b2ef6,
24'h3b2ef6,
24'h3b2ef6,
24'h4e4dff,
24'h4e4dff,
24'h4e47ff,
24'h4e47ff,
24'h4e47ff,
24'h4a3dee,
24'h4a3dee,
24'h4735ff,
24'h4735ff,
24'h4735ff,
24'h4235fd,
24'h4235fd,
24'h4237fc,
24'h4237fc,
24'h4237fc,
24'h4338fd,
24'h4338fd,
24'h4336ff,
24'h4336ff,
24'h4336ff,
24'h493aff,
24'h493aff,
24'h4e43ff,
24'h4e43ff,
24'h4e43ff,
24'h4d47ff,
24'h4d47ff,
24'h4540fd,
24'h4540fd,
24'h4540fd,
24'h4539fe,
24'h4539fe,
24'h422ffa,
24'h422ffa,
24'h422ffa,
24'h463aff,
24'h463aff,
24'h3b2ef6,
24'h3b2ef6,
24'h3b2ef6,
24'h4e4dff,
24'h4e4dff,
24'h4e47ff,
24'h4e47ff,
24'h4e47ff,
24'h4a3dee,
24'h4a3dee,
24'h4735ff,
24'h4735ff,
24'h4735ff,
24'h4235fd,
24'h4235fd,
24'h4237fc,
24'h4237fc,
24'h4237fc,
24'h4338fd,
24'h4338fd,
24'h4336ff,
24'h4336ff,
24'h4336ff,
24'h493aff,
24'h493aff,
24'h4e43ff,
24'h4e43ff,
24'h4e43ff,
24'h4d47ff,
24'h4d47ff,
24'h4540fd,
24'h4540fd,
24'h4540fd,
24'h4539fe,
24'h4539fe,
24'h422ffa,
24'h422ffa,
24'h422ffa,
24'h4933ff,
24'h4933ff,
24'h3a44ff,
24'h3a44ff,
24'h3a44ff,
24'h4042ff,
24'h4042ff,
24'h4b3aff,
24'h4b3aff,
24'h4b3aff,
24'h4636f8,
24'h4636f8,
24'h4737ff,
24'h4737ff,
24'h4737ff,
24'h4437ff,
24'h4437ff,
24'h4138ff,
24'h4138ff,
24'h4138ff,
24'h4037ff,
24'h4037ff,
24'h3e32ff,
24'h3e32ff,
24'h3e32ff,
24'h4032ff,
24'h4032ff,
24'h3e35ff,
24'h3e35ff,
24'h3e35ff,
24'h3733f8,
24'h3733f8,
24'h3c35f4,
24'h3c35f4,
24'h3c35f4,
24'h3e31f9,
24'h3e31f9,
24'h4b35ff,
24'h4b35ff,
24'h4b35ff,
24'h4933ff,
24'h4933ff,
24'h3a44ff,
24'h3a44ff,
24'h3a44ff,
24'h4042ff,
24'h4042ff,
24'h4b3aff,
24'h4b3aff,
24'h4b3aff,
24'h4636f8,
24'h4636f8,
24'h4737ff,
24'h4737ff,
24'h4737ff,
24'h4437ff,
24'h4437ff,
24'h4138ff,
24'h4138ff,
24'h4138ff,
24'h4037ff,
24'h4037ff,
24'h3e32ff,
24'h3e32ff,
24'h3e32ff,
24'h4032ff,
24'h4032ff,
24'h3e35ff,
24'h3e35ff,
24'h3e35ff,
24'h3733f8,
24'h3733f8,
24'h3c35f4,
24'h3c35f4,
24'h3c35f4,
24'h3e31f9,
24'h3e31f9,
24'h4b35ff,
24'h4b35ff,
24'h4b35ff,
24'h3f2fff,
24'h3f2fff,
24'h393efb,
24'h393efb,
24'h393efb,
24'h4130f1,
24'h4130f1,
24'h4b32ff,
24'h4b32ff,
24'h4b32ff,
24'h3a30ff,
24'h3a30ff,
24'h4134f5,
24'h4134f5,
24'h4134f5,
24'h483ffd,
24'h483ffd,
24'h504aff,
24'h504aff,
24'h504aff,
24'h504aff,
24'h504aff,
24'h4a41ff,
24'h4a41ff,
24'h4a41ff,
24'h4b3fff,
24'h4b3fff,
24'h4e47ff,
24'h4e47ff,
24'h4e47ff,
24'h4d4bff,
24'h4d4bff,
24'h3e33f8,
24'h3e33f8,
24'h3e33f8,
24'h4b3cff,
24'h4b3cff,
24'h4630fe,
24'h4630fe,
24'h4630fe,
24'h3f2fff,
24'h3f2fff,
24'h393efb,
24'h393efb,
24'h393efb,
24'h4130f1,
24'h4130f1,
24'h4b32ff,
24'h4b32ff,
24'h4b32ff,
24'h3a30ff,
24'h3a30ff,
24'h4134f5,
24'h4134f5,
24'h4134f5,
24'h483ffd,
24'h483ffd,
24'h504aff,
24'h504aff,
24'h504aff,
24'h504aff,
24'h504aff,
24'h4a41ff,
24'h4a41ff,
24'h4a41ff,
24'h4b3fff,
24'h4b3fff,
24'h4e47ff,
24'h4e47ff,
24'h4e47ff,
24'h4d4bff,
24'h4d4bff,
24'h3e33f8,
24'h3e33f8,
24'h3e33f8,
24'h4b3cff,
24'h4b3cff,
24'h4630fe,
24'h4630fe,
24'h4630fe,
24'h3f2fff,
24'h3f2fff,
24'h393efb,
24'h393efb,
24'h393efb,
24'h4130f1,
24'h4130f1,
24'h4b32ff,
24'h4b32ff,
24'h4b32ff,
24'h3a30ff,
24'h3a30ff,
24'h4134f5,
24'h4134f5,
24'h4134f5,
24'h483ffd,
24'h483ffd,
24'h504aff,
24'h504aff,
24'h504aff,
24'h504aff,
24'h504aff,
24'h4a41ff,
24'h4a41ff,
24'h4a41ff,
24'h4b3fff,
24'h4b3fff,
24'h4e47ff,
24'h4e47ff,
24'h4e47ff,
24'h4d4bff,
24'h4d4bff,
24'h3e33f8,
24'h3e33f8,
24'h3e33f8,
24'h4b3cff,
24'h4b3cff,
24'h4630fe,
24'h4630fe,
24'h4630fe,
24'h4832ff,
24'h4832ff,
24'h4333f5,
24'h4333f5,
24'h4333f5,
24'h5746ff,
24'h5746ff,
24'h4e45ff,
24'h4e45ff,
24'h4e45ff,
24'h4c49ff,
24'h4c49ff,
24'h4438fd,
24'h4438fd,
24'h4438fd,
24'h463ffe,
24'h463ffe,
24'h4a45ff,
24'h4a45ff,
24'h4a45ff,
24'h4841ff,
24'h4841ff,
24'h4337fc,
24'h4337fc,
24'h4337fc,
24'h4336fe,
24'h4336fe,
24'h4439fe,
24'h4439fe,
24'h4439fe,
24'h413afb,
24'h413afb,
24'h4338ff,
24'h4338ff,
24'h4338ff,
24'h4334ff,
24'h4334ff,
24'h452dfc,
24'h452dfc,
24'h452dfc,
24'h4832ff,
24'h4832ff,
24'h4333f5,
24'h4333f5,
24'h4333f5,
24'h5746ff,
24'h5746ff,
24'h4e45ff,
24'h4e45ff,
24'h4e45ff,
24'h4c49ff,
24'h4c49ff,
24'h4438fd,
24'h4438fd,
24'h4438fd,
24'h463ffe,
24'h463ffe,
24'h4a45ff,
24'h4a45ff,
24'h4a45ff,
24'h4841ff,
24'h4841ff,
24'h4337fc,
24'h4337fc,
24'h4337fc,
24'h4336fe,
24'h4336fe,
24'h4439fe,
24'h4439fe,
24'h4439fe,
24'h413afb,
24'h413afb,
24'h4338ff,
24'h4338ff,
24'h4338ff,
24'h4334ff,
24'h4334ff,
24'h452dfc,
24'h452dfc,
24'h452dfc,
24'h412aeb,
24'h412aeb,
24'h473aff,
24'h473aff,
24'h473aff,
24'h3c39ff,
24'h3c39ff,
24'h383dfa,
24'h383dfa,
24'h383dfa,
24'h3d33f5,
24'h3d33f5,
24'h4135ff,
24'h4135ff,
24'h4135ff,
24'h3d34fc,
24'h3d34fc,
24'h3c36fb,
24'h3c36fb,
24'h3c36fb,
24'h3c33fb,
24'h3c33fb,
24'h3f31ff,
24'h3f31ff,
24'h3f31ff,
24'h4835ff,
24'h4835ff,
24'h4636ff,
24'h4636ff,
24'h4636ff,
24'h3e32ff,
24'h3e32ff,
24'h3f32fb,
24'h3f32fb,
24'h3f32fb,
24'h4634ff,
24'h4634ff,
24'h4830ff,
24'h4830ff,
24'h4830ff,
24'h412aeb,
24'h412aeb,
24'h473aff,
24'h473aff,
24'h473aff,
24'h3c39ff,
24'h3c39ff,
24'h383dfa,
24'h383dfa,
24'h383dfa,
24'h3d33f5,
24'h3d33f5,
24'h4135ff,
24'h4135ff,
24'h4135ff,
24'h3d34fc,
24'h3d34fc,
24'h3c36fb,
24'h3c36fb,
24'h3c36fb,
24'h3c33fb,
24'h3c33fb,
24'h3f31ff,
24'h3f31ff,
24'h3f31ff,
24'h4835ff,
24'h4835ff,
24'h4636ff,
24'h4636ff,
24'h4636ff,
24'h3e32ff,
24'h3e32ff,
24'h3f32fb,
24'h3f32fb,
24'h3f32fb,
24'h4634ff,
24'h4634ff,
24'h4830ff,
24'h4830ff,
24'h4830ff,
24'h412aeb,
24'h412aeb,
24'h473aff,
24'h473aff,
24'h473aff,
24'h3c39ff,
24'h3c39ff,
24'h383dfa,
24'h383dfa,
24'h383dfa,
24'h3d33f5,
24'h3d33f5,
24'h4135ff,
24'h4135ff,
24'h4135ff,
24'h3d34fc,
24'h3d34fc,
24'h3c36fb,
24'h3c36fb,
24'h3c36fb,
24'h3c33fb,
24'h3c33fb,
24'h3f31ff,
24'h3f31ff,
24'h3f31ff,
24'h4835ff,
24'h4835ff,
24'h4636ff,
24'h4636ff,
24'h4636ff,
24'h3e32ff,
24'h3e32ff,
24'h3f32fb,
24'h3f32fb,
24'h3f32fb,
24'h4634ff,
24'h4634ff,
24'h4830ff,
24'h4830ff,
24'h4830ff,
24'h4d48fc,
24'h4d48fc,
24'h4048ff,
24'h4048ff,
24'h4048ff,
24'h4646ff,
24'h4646ff,
24'h4543fb,
24'h4543fb,
24'h4543fb,
24'h5347fe,
24'h5347fe,
24'h4e45ff,
24'h4e45ff,
24'h4e45ff,
24'h4c46ff,
24'h4c46ff,
24'h4a45ff,
24'h4a45ff,
24'h4a45ff,
24'h453efc,
24'h453efc,
24'h4335fb,
24'h4335fb,
24'h4335fb,
24'h4736ff,
24'h4736ff,
24'h4837ff,
24'h4837ff,
24'h4837ff,
24'h4034f9,
24'h4034f9,
24'h4033fe,
24'h4033fe,
24'h4033fe,
24'h4331ff,
24'h4331ff,
24'h4d35ff,
24'h4d35ff,
24'h4d35ff,
24'h4d48fc,
24'h4d48fc,
24'h4048ff,
24'h4048ff,
24'h4048ff,
24'h4646ff,
24'h4646ff,
24'h4543fb,
24'h4543fb,
24'h4543fb,
24'h5347fe,
24'h5347fe,
24'h4e45ff,
24'h4e45ff,
24'h4e45ff,
24'h4c46ff,
24'h4c46ff,
24'h4a45ff,
24'h4a45ff,
24'h4a45ff,
24'h453efc,
24'h453efc,
24'h4335fb,
24'h4335fb,
24'h4335fb,
24'h4736ff,
24'h4736ff,
24'h4837ff,
24'h4837ff,
24'h4837ff,
24'h4034f9,
24'h4034f9,
24'h4033fe,
24'h4033fe,
24'h4033fe,
24'h4331ff,
24'h4331ff,
24'h4d35ff,
24'h4d35ff,
24'h4d35ff,
24'h3f32ff,
24'h3f32ff,
24'h452ffb,
24'h452ffb,
24'h452ffb,
24'h4d2cff,
24'h4d2cff,
24'h4436ff,
24'h4436ff,
24'h4436ff,
24'h3f32fa,
24'h3f32fa,
24'h403bf9,
24'h403bf9,
24'h403bf9,
24'h433efc,
24'h433efc,
24'h4742ff,
24'h4742ff,
24'h4742ff,
24'h4b46ff,
24'h4b46ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4c47ff,
24'h4c47ff,
24'h4c47ff,
24'h4a45ff,
24'h4a45ff,
24'h433dff,
24'h433dff,
24'h433dff,
24'h4034ff,
24'h4034ff,
24'h4737f8,
24'h4737f8,
24'h4737f8,
24'h3f32ff,
24'h3f32ff,
24'h452ffb,
24'h452ffb,
24'h452ffb,
24'h4d2cff,
24'h4d2cff,
24'h4436ff,
24'h4436ff,
24'h4436ff,
24'h3f32fa,
24'h3f32fa,
24'h403bf9,
24'h403bf9,
24'h403bf9,
24'h433efc,
24'h433efc,
24'h4742ff,
24'h4742ff,
24'h4742ff,
24'h4b46ff,
24'h4b46ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4c47ff,
24'h4c47ff,
24'h4c47ff,
24'h4a45ff,
24'h4a45ff,
24'h433dff,
24'h433dff,
24'h433dff,
24'h4034ff,
24'h4034ff,
24'h4737f8,
24'h4737f8,
24'h4737f8,
24'h3f32ff,
24'h3f32ff,
24'h452ffb,
24'h452ffb,
24'h452ffb,
24'h4d2cff,
24'h4d2cff,
24'h4436ff,
24'h4436ff,
24'h4436ff,
24'h3f32fa,
24'h3f32fa,
24'h403bf9,
24'h403bf9,
24'h403bf9,
24'h433efc,
24'h433efc,
24'h4742ff,
24'h4742ff,
24'h4742ff,
24'h4b46ff,
24'h4b46ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4d48ff,
24'h4c47ff,
24'h4c47ff,
24'h4c47ff,
24'h4a45ff,
24'h4a45ff,
24'h433dff,
24'h433dff,
24'h433dff,
24'h4034ff,
24'h4034ff,
24'h4737f8,
24'h4737f8,
24'h4737f8,
24'h363fff,
24'h363fff,
24'h3943f1,
24'h3943f1,
24'h3943f1,
24'h4f40fa,
24'h4f40fa,
24'h4c49ff,
24'h4c49ff,
24'h4c49ff,
24'h4448ff,
24'h4448ff,
24'h493cff,
24'h493cff,
24'h493cff,
24'h473aff,
24'h473aff,
24'h4336fe,
24'h4336fe,
24'h4336fe,
24'h4033fb,
24'h4033fb,
24'h3f32fa,
24'h3f32fa,
24'h3f32fa,
24'h4034f9,
24'h4034f9,
24'h4337fc,
24'h4337fc,
24'h4337fc,
24'h4438fd,
24'h4438fd,
24'h3d32f9,
24'h3d32f9,
24'h3d32f9,
24'h5342ff,
24'h5342ff,
24'h5440ff,
24'h5440ff,
24'h5440ff,
24'h363fff,
24'h363fff,
24'h3943f1,
24'h3943f1,
24'h3943f1,
24'h4f40fa,
24'h4f40fa,
24'h4c49ff,
24'h4c49ff,
24'h4c49ff,
24'h4448ff,
24'h4448ff,
24'h493cff,
24'h493cff,
24'h493cff,
24'h473aff,
24'h473aff,
24'h4336fe,
24'h4336fe,
24'h4336fe,
24'h4033fb,
24'h4033fb,
24'h3f32fa,
24'h3f32fa,
24'h3f32fa,
24'h4034f9,
24'h4034f9,
24'h4337fc,
24'h4337fc,
24'h4337fc,
24'h4438fd,
24'h4438fd,
24'h3d32f9,
24'h3d32f9,
24'h3d32f9,
24'h5342ff,
24'h5342ff,
24'h5440ff,
24'h5440ff,
24'h5440ff,
24'h472bf9,
24'h472bf9,
24'h462bff,
24'h462bff,
24'h462bff,
24'h4c2eff,
24'h4c2eff,
24'h4538ff,
24'h4538ff,
24'h4538ff,
24'h4134ff,
24'h4134ff,
24'h4c39ff,
24'h4c39ff,
24'h4c39ff,
24'h4a37ff,
24'h4a37ff,
24'h4835ff,
24'h4835ff,
24'h4835ff,
24'h4532fd,
24'h4532fd,
24'h4431fc,
24'h4431fc,
24'h4431fc,
24'h4532fd,
24'h4532fd,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4433fd,
24'h4433fd,
24'h4433fd,
24'h4a33ff,
24'h4a33ff,
24'h4834e2,
24'h4834e2,
24'h4834e2,
24'h472bf9,
24'h472bf9,
24'h462bff,
24'h462bff,
24'h462bff,
24'h4c2eff,
24'h4c2eff,
24'h4538ff,
24'h4538ff,
24'h4538ff,
24'h4134ff,
24'h4134ff,
24'h4c39ff,
24'h4c39ff,
24'h4c39ff,
24'h4a37ff,
24'h4a37ff,
24'h4835ff,
24'h4835ff,
24'h4835ff,
24'h4532fd,
24'h4532fd,
24'h4431fc,
24'h4431fc,
24'h4431fc,
24'h4532fd,
24'h4532fd,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4433fd,
24'h4433fd,
24'h4433fd,
24'h4a33ff,
24'h4a33ff,
24'h4834e2,
24'h4834e2,
24'h4834e2,
24'h472bf9,
24'h472bf9,
24'h462bff,
24'h462bff,
24'h462bff,
24'h4c2eff,
24'h4c2eff,
24'h4538ff,
24'h4538ff,
24'h4538ff,
24'h4134ff,
24'h4134ff,
24'h4c39ff,
24'h4c39ff,
24'h4c39ff,
24'h4a37ff,
24'h4a37ff,
24'h4835ff,
24'h4835ff,
24'h4835ff,
24'h4532fd,
24'h4532fd,
24'h4431fc,
24'h4431fc,
24'h4431fc,
24'h4532fd,
24'h4532fd,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4633ff,
24'h4433fd,
24'h4433fd,
24'h4433fd,
24'h4a33ff,
24'h4a33ff,
24'h4834e2,
24'h4834e2,
24'h4834e2
};
parameter bit [23:0] rom_chest[1599:0]
='{24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'ha47227,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17,
24'h211d17
};
parameter bit [23:0] rom_wooden_planks[1599:0]
='{24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'hbc9862,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a
};
always_comb
begin
 if(rely<40&relx<40)	
 begin
	case(id)

	4'd1:
		rgb= rom_bedrock[rely*40+relx];
	4'd2:
		rgb= rom_wood [rely*40+relx];
	4'd3:
		rgb= rom_stone [rely*40+relx];
	4'd4:
		rgb= rom_dirt [rely*40+relx];
	4'd5:
		rgb= rom_diamond_ore [rely*40+relx];
	4'd6:
		rgb= rom_furnace [rely*40+relx];
	4'd7:
		rgb= rom_gold_ore [rely*40+relx];	
	4'd8:
		rgb= rom_grass [rely*40+relx];
	4'd9:
		rgb= rom_iron_ore [rely*40+relx];
	4'd10:
		rgb= rom_leaves [rely*40+relx];
	4'd11:
		rgb= rom_coal_ore [rely*40+relx];
	4'd12:
		rgb= rom_crafting_table [rely*40+relx];
	4'd13:
		rgb= rom_water [rely*40+relx];
	4'd14:
		rgb= rom_chest [rely*40+relx];
	4'd15:
		rgb= rom_wooden_planks [rely*40+relx];
	default:
		rgb=0;
	endcase
	
 end
 else
 
 rgb=24'b0;
 
end

always_comb
begin
	if((steve_relx!=6'b0)&(steve_rely!=6'b0))
	begin
		steve_rgb=rom_steve[(79-steve_rely)*40+steve_relx];
	end
	
	else
		steve_rgb=24'hd2e6ff;
end







endmodule