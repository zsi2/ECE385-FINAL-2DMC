module false_map

(

	input logic [9:0] corner_x,corner_y, // lefttop corner of buffer
	
	output logic [63:0] row_0,row_1,row_2,row_3,row_4,row_5,row_6,row_7,row_8,row_9,row_10,row_11,
	
	input logic [9:0] changex,changey,
	
	input logic [1:0]operation,
	input logic Clk,Reset_h,
	
	input logic [3:0] push_id


);

/*parameter bit [31:0] map_tile0 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h80000000,
32'hC8000000,
32'hCC888000,
32'hCBCCC888,
32'hCBBCCCCC,
32'hBBBCCBCC,
32'hBBBBCBBC,
32'hBBBBBBBC,
32'hBBBBBBBC,
32'hBBBBBBBB,
32'hB9BBBB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB3BB,
32'hBB93BBB9,
32'hBBBBBBB3,
32'hBBBBBBB3,
32'hB7BBBBBB,
32'h7BB9BBBB,
32'hBBBBBBBB,
32'hBBB7BBBB,
32'hBBBBBBBB,
32'hBBBBBB37,
32'hBBBB7BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hBBBBBBB7,
32'hBBB3BBBB,
32'hBBBBB9B5,
32'hBB3BBB33,
32'hBBBBBB77,
32'hBBBB9BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hB3BBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB7BB7BB,
32'hBBB9BBBB,
32'hBB5BBB9B,
32'h9BBB5BBB,
32'hBBB9BBBB,
32'h11111111
};
parameter bit [31:0] map_tile1 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h0000000A,
32'h000000AA,
32'h00000AAA,
32'h08880000,
32'h0CCC0000,
32'h8CCC8800,
32'hCCCCCC88,
32'hCBCCBBCC,
32'hCBBBBBCC,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB9BBBBBB,
32'hBBBBBBBB,
32'hBBB3BBBB,
32'hBB39BBBB,
32'hBBBBBBBB,
32'h3BBBBBB9,
32'hBBBBBBBB,
32'hBBBBBB3B,
32'hBBBB73BB,
32'hB3BBBBBB,
32'hBBBBBBBB,
32'hBBBBBB3B,
32'hBBBBBBBB,
32'hBBB39BBB,
32'hBB9BBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB33B,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hBBBB9BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB9BBBBB,
32'hBBB7B9BB,
32'hBBBBBBBB,
32'hB37BBBBB,
32'hBBBBBBBB,
32'hBBB7BB7B,
32'hBBBB53BB,
32'hBBBB9BBB,
32'hBB3BBBBB,
32'h5BB9BBBB,
32'hBB7BBBBB,
32'hBBB9BBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB9BBBB,
32'hBBBBBBB7,
32'hBBBB3BBB,
32'h11111111
};
parameter bit [31:0] map_tile2 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'hA0000000,
32'hAA000000,
32'hEAA00000,
32'hEAAA0000,
32'hE0000000,
32'hE0000088,
32'hE08000CC,
32'h88C088CC,
32'hCCC8CCBC,
32'hBCBCCCBC,
32'hBBBBBCBC,
32'hBBBBBB9B,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'hBBBB9BBB,
32'hBBBBBB3B,
32'hBBB799BB,
32'hBBBBB7BB,
32'hBBBBBBBB,
32'h3BBBB3BB,
32'hBBBBBBBB,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB7BBBB,
32'hBBBBBB3B,
32'hBBBBB3BB,
32'h7BBBBB9B,
32'hBBBBBBBB,
32'hBBBBBB9B,
32'hBBBBBB9B,
32'hB7BB7BBB,
32'hBBBBBBBB,
32'hB9BBBBBB,
32'hBBB9BBB3,
32'hBBBBBBBB,
32'hBBBBBB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB3BBBB9,
32'hBBBBBB5B,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'hBBBB5BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h3BB9BBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB7BB,
32'hBB9BBBBB,
32'hBBBBBBB3,
32'hB3BBBBBB,
32'hBBBBBBBB,
32'h11111111
};
parameter bit [31:0] map_tile3 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000088,
32'h008008CC,
32'h88C88CCB,
32'hCCCCCCBB,
32'hCCCCCBBB,
32'hCCCCCBBB,
32'hBBCCCBBB,
32'hBBBCCBB3,
32'hBB9BBBBB,
32'hB9BBBBBB,
32'hBBBBBBB9,
32'hBBBBBBBB,
32'h7BBB3BBB,
32'hBBBBBBBB,
32'h7BBBBBBB,
32'hBB3BB3BB,
32'hBB3BBBBB,
32'hBB3BBBBB,
32'h9B3BB7BB,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'hBBBBBBBB,
32'h373BBBBB,
32'hB3BBB33B,
32'hB7BBB3BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB3BBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB77B9BBB,
32'hBBBBB3BB,
32'hBB9BBB3B,
32'hB3BBBBBB,
32'h7BBB33BB,
32'hBBB33BBB,
32'hB3BBBB9B,
32'hBBBBB3BB,
32'hBBBBBBBB,
32'hB3BBBBBB,
32'hBBBBBBBB,
32'hB9BBBBB3,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hB5BBBBBB,
32'h9BBBBBBB,
32'hBB9BBBBB,
32'hBB33BBBB,
32'hB3B5BBBB,
32'hBBBBBBBB,
32'hBBBBB7BB,
32'h11111111
};
parameter bit [31:0] map_tile4 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000088,
32'h808888CC,
32'hC8CCCCCC,
32'hCCCCCBBC,
32'hBCCCCBBC,
32'hBCBCBBBB,
32'hBCBCBBBB,
32'hBCBBBBBB,
32'hBBBBBBBB,
32'hBBB9BBBB,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBB7BBB,
32'hBBBBBBBB,
32'hBBBB3BBB,
32'hBBBBBB9B,
32'h7BBBB3BB,
32'h9BBBBBBB,
32'hBBBBBBBB,
32'hBBB9BBBB,
32'h9BBBBBBB,
32'hBBBBBBBB,
32'h3BB3BBBB,
32'hB9BBB3B9,
32'hBBBBBBBB,
32'hBB7BBB3B,
32'h3B3BBB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBB7B,
32'hBBBBBBBB,
32'hBB9BBBBB,
32'h9BBBBBBB,
32'hBB9BBBBB,
32'hBBBB99BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h5BBBBB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBB77,
32'hBBBB35B7,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB5BBB7B,
32'hBBB7BBB3,
32'hBBB5BBBB,
32'h11111111
};
parameter bit [31:0] map_tile5 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h0000000A,
32'h000000AA,
32'h00000AAE,
32'h0000AAAE,
32'h0000000E,
32'h0888000E,
32'h8CCC880E,
32'hCCCBCC88,
32'hBBCBCCCC,
32'hBBBBBCCC,
32'hBBBBBBBC,
32'hBBB9BBBC,
32'hB9BBBBBB,
32'hBB9BBBB3,
32'hBBB9BBBB,
32'hBBBB3B39,
32'hBBBBBBBB,
32'hBBBBBB93,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'hBBBB3BBB,
32'hBBB9BBBB,
32'hBBB3BBBB,
32'hB9BBBBBB,
32'hBBBB3B3B,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBB9BBB,
32'hBBBBB7B3,
32'hBB9BBB3B,
32'h3BBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBB3B,
32'h3BBBBBBB,
32'h3BBBBB3B,
32'hBBBBBB93,
32'hB3BBBBBB,
32'hBBBB9BBB,
32'hBBBBBBB9,
32'hBBBB3BBB,
32'hBBBBBBBB,
32'hBBBBBB3B,
32'hB7BBBB5B,
32'hB3BBBBBB,
32'hBBB9BBBB,
32'hB9BBBBBB,
32'hBBBB3BBB,
32'hBBBBBBBB,
32'hBBBBB93B,
32'h3BBBBBBB,
32'hBB3BBBBB,
32'hBBB5BBB3,
32'h3BBBBBBB,
32'hBBBBBBBB,
32'hBB3BBB33,
32'hB7BBB3BB,
32'h11111111
};
parameter bit [31:0] map_tile6 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'hA0000000,
32'hAA000088,
32'hAAA000CC,
32'h000008CC,
32'h00008CCC,
32'h0008CCCB,
32'h800CCCCB,
32'hC88CCCBB,
32'hBCCCBCBB,
32'hBCCCBBBB,
32'hBCCBBBBB,
32'hBBCBBBBB,
32'hBBBBBBBB,
32'h93BBBBBB,
32'hBBBBBBBB,
32'h3BBB3B3B,
32'hBBBB3BBB,
32'h3BBB3BBB,
32'hBBBB9B33,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBB3B,
32'hBBBBBBBB,
32'hBBBBBBB9,
32'hB3B9B7BB,
32'hBBB9B93B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB7B7B3BB,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'hBBBBBBBB,
32'hB39BBBBB,
32'hBB9BBBBB,
32'hB7BBBBBB,
32'h7BB9BBBB,
32'h3BBBBBBB,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBB9BBB,
32'hBBBBB3BB,
32'hBBBBBB7B,
32'h99BBBB3B,
32'hBBBBBB3B,
32'hBB5BBBBB,
32'hBBBBBB5B,
32'h5BBBBBBB,
32'hBBBBB3BB,
32'hBBBBBB3B,
32'hB5BBBBBB,
32'hBBBB5BBB,
32'hBBBBBBBB,
32'h5BBBBBBB,
32'h11111111
};
parameter bit [31:0] map_tile7 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h000A0000,
32'h00AAA000,
32'h0AAEAA00,
32'hAAAEAAA0,
32'h000E0000,
32'h000E0000,
32'h000E0088,
32'h888888CC,
32'hCCCCCCCC,
32'hCCCBCBCC,
32'hCCBBCBCB,
32'hCCBBBBCB,
32'hCCBBBBBB,
32'hBBBBB9B3,
32'hBBBBBBBB,
32'h3BBB3B3B,
32'hBBBBBBBB,
32'hBBBBB39B,
32'hB3BBBB3B,
32'h3B9BB9B9,
32'hBB9BBB3B,
32'hBBB3BBBB,
32'hBB3B3BBB,
32'hBBB3BBB9,
32'hBBBBB3BB,
32'hBBBB3BBB,
32'hBBB3BBBB,
32'hB7BBBBBB,
32'hBBBB7BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB3BBBBBB,
32'hB9BBBBB9,
32'hBB3BB7BB,
32'hBB3BB3BB,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hBBBBBB7B,
32'hBB3BBBB9,
32'hBBBBBBBB,
32'hBBBBB9BB,
32'hBBBBBB3B,
32'hBB9B3BBB,
32'hBB7BBBBB,
32'hBB3BBBBB,
32'hBBBB7BBB,
32'hBB3BBBBB,
32'hB9BBBBBB,
32'hBBBBBBBB,
32'hBBBBBBB9,
32'hBBB9B7BB,
32'hBBBB7B3B,
32'hBBBB3BBB,
32'hBBBBBBBB,
32'h7BBBBBBB,
32'hBBBBBBBB,
32'h37B39BBB,
32'hBBBBBBBB,
32'hBBB7B37B,
32'hBBBBB3BB,
32'hBBBBBBB5,
32'hBBBBBBBB,
32'h11111111
};
parameter bit [31:0] map_tile8 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h88808880,
32'hCCC8CCC0,
32'hCCCCCCC8,
32'hCCCCBCCC,
32'hBCBCBCCC,
32'hBBBBBBCC,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB93BBB,
32'hB3BBBBBB,
32'hB3BBBBB3,
32'hBBBBBBB9,
32'hBBB3BB3B,
32'hBBBBBBBB,
32'hB3BBBBBB,
32'hBBBB33BB,
32'hB3BBB3B3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB3B3BB,
32'hBBBBBBB7,
32'hBBBBBBB9,
32'hB3BB33BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h3BBBBBB9,
32'hB7B7BBBB,
32'hBBB7BBBB,
32'hB7BBBBBB,
32'hBBBBBBB3,
32'hBB9B9BBB,
32'hBB9BB9BB,
32'h3BBBBBBB,
32'hBBBBB7BB,
32'hBBBBBBBB,
32'hBBBBBBB9,
32'h9BBBBBBB,
32'hB7BBB9BB,
32'hBBBBBB3B,
32'hBBBBBB9B,
32'hBBBBBBB5,
32'hBB3BBBBB,
32'hBB7BBBBB,
32'hBBBBBBBB,
32'h3BBBBBB9,
32'hB3BB7BBB,
32'hBBBB3BBB,
32'hBBB9BBBB,
32'hB9BBBBBB,
32'h3BBBBBBB,
32'hBBBBBBBB,
32'h93BBBBBB,
32'hBBB5BBBB,
32'h7BBBBBBB,
32'hBBBB5BBB,
32'hBBB3BBBB,
32'h9BBBB5BB,
32'hBBBB3BBB,
32'h11111111
};
parameter bit [31:0] map_tile9 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000088,
32'h000088CC,
32'h0080CCCC,
32'h88C8CCCC,
32'hCCCCCCCC,
32'hCCBBCCBB,
32'hBCBBBBB3,
32'hBCBBBBBB,
32'hBBBB3BBB,
32'hBBBB9B3B,
32'hBBB99BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB3BB,
32'hBBBBBBBB,
32'hBBBBBB9B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBB9,
32'h7BBBBBBB,
32'hB9BBBBBB,
32'hB3BB3B93,
32'hBBBBBBBB,
32'hB3BBBBB9,
32'hBBBBB33B,
32'hBBBBB93B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB7BBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB9BB7B9,
32'h7BBBBBBB,
32'hBBBBBBB9,
32'hBBBBBBB3,
32'hBB3BBBBB,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBB9B7B,
32'hBBBB5BB3,
32'hBBBBBB3B,
32'h53BBBBBB,
32'hBBBBBBBB,
32'hBBBB5BBB,
32'hBBBB97BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB9BBB9B3,
32'hBBBBBBB3,
32'hBBBBB3B3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBB7B,
32'hBBBBBB5B,
32'h99BB7BB3,
32'h9BBBBBBB,
32'hBB3BBBBB,
32'h11111111
};
parameter bit [31:0] map_tile10 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h0000000A,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00080000,
32'h888C8888,
32'hCCCCCCCC,
32'hCCBCCCCC,
32'hCCBCCCBC,
32'hCCBBCCBC,
32'hBBBBBCBC,
32'hBB3BBB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB3BBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB9BB,
32'h33BBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBB3BBB,
32'hBBBBBBBB,
32'hBBBBBB3B,
32'hBBBBBBBB,
32'h79BBBBBB,
32'hBBB9BB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBB3BBB,
32'h33BBBBBB,
32'h9BBBBBBB,
32'hBBBBBBBB,
32'hBB9BBBBB,
32'hBB7BBBBB,
32'hBBBBB3BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h3B3BBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB3BBBB,
32'hBB93BBBB,
32'hBBBBBBBB,
32'hBBBBBB9B,
32'h7BBBBBB9,
32'hBBB3B9BB,
32'hBBBB3BB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBB5B,
32'hBBB9BBB3,
32'hBBB9BBBB,
32'hB3BBB357,
32'hBB9BBBBB,
32'hBBBBB35B,
32'hBB7BBBBB,
32'hBBBBBBBB,
32'h5BBBBBBB,
32'hBBBBBBBB,
32'h11111111
};
parameter bit [31:0] map_tile11 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00A00000,
32'h0AAA0000,
32'hAAEAA000,
32'hAAEAAA00,
32'h00E00000,
32'h00E00000,
32'h00E00000,
32'h88800000,
32'hCCC80000,
32'hCCCC8000,
32'hCCCCC888,
32'hBBBCCCCC,
32'hBBBCCBCC,
32'hBBBBBBCC,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hBBB3BBBB,
32'hBB3BBBBB,
32'hBBBBBBB9,
32'hBBBBB9BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h93BBB33B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB3BB,
32'hBBBBBBBB,
32'hBBBBBBB9,
32'h79BBBBBB,
32'hBBBBBBBB,
32'hBBBB33BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB9BBB9B,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBB3BBB,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hBBB9BBBB,
32'hBBB3BB37,
32'hBB7BBB73,
32'hBBBBBB3B,
32'hB3BBBBBB,
32'hBBBBBBB7,
32'hB3BB7BBB,
32'hB9BB9BBB,
32'hBBBBBBBB,
32'hBB3BB3BB,
32'hBBB5BBBB,
32'hBBB9BBBB,
32'hBBBB3BBB,
32'hBBBBBB9B,
32'hBB7BBBBB,
32'hBBBBB9BB,
32'hBBBBB7BB,
32'hBBBBB9BB,
32'hBBBBBB7B,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'h3BBB7BBB,
32'h11111111
};
parameter bit [31:0] map_tile12[99:0] ='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00008000,
32'h8888C888,
32'hCCCCCCCC,
32'hCCBCCCCC,
32'hBCBCCCBC,
32'hBCBCCBBC,
32'hBBBBBBBC,
32'hBBBBBBBB,
32'hBBBBB9BB,
32'hBBBBBBBB,
32'hBB3BB3B9,
32'hBBBBBBBB,
32'hBBB3BBBB,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'hBBBBBBBB,
32'hBB9BBBBB,
32'hBBBBB3B9,
32'hBB3BBBBB,
32'hBBBBB3BB,
32'hBBBBBBBB,
32'hBB99BBBB,
32'hB3BBBBBB,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB3BBBB,
32'hBBBBB7B3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'hB3BBBBBB,
32'hBB7BBBBB,
32'hBBBB9B7B,
32'h9BBBBBB3,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'h9BBB9BB3,
32'hBBBBBBB7,
32'hBBBBBBBB,
32'hB7BB3BBB,
32'hBBBBBB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h3BBBBBB7,
32'hBBB9BB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBB3BBB,
32'hBBBBB5B3,
32'h9BBBBBB3,
32'h9BBBBB5B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB39B,
32'hB3BBBBBB,
32'h3BB7BBBB,
32'hBBBBBBBB,
32'h11111111
};
parameter bit [31:0] map_tile13 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000888,
32'h88888CCC,
32'hCCCCCCCB,
32'hCCCBCCCB,
32'hBCCBCCBB,
32'hBBCBCCBB,
32'hBBCBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB9BBBBBB,
32'hBBBBBBB9,
32'h3BBBBBBB,
32'h3BBBBB3B,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hBBBBBBB9,
32'h3BBBBBB3,
32'hBBBBBBBB,
32'h3BBBBBBB,
32'hBBB9B3BB,
32'hBBBBBBBB,
32'hB3B9BBBB,
32'h3BBB9BBB,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hBB9B3BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB9BBBBB,
32'hBBB3BB9B,
32'hBBB3BBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB33BB93B,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hB7BBBBBB,
32'hBBBBB3BB,
32'hBBBBBBBB,
32'h3BBBBB9B,
32'hBBBBB3BB,
32'hBBBBBBBB,
32'hBBBB9B3B,
32'hBBBBBBB5,
32'hB3BBBBBB,
32'hB3BB7BB9,
32'hBBB3BBBB,
32'hBBBBBBBB,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'h5BBBB3BB,
32'hBBBBBBBB,
32'h9BBBBBB7,
32'hB3BBBBB9,
32'hB3BB5BB7,
32'hBBB7B35B,
32'hBBBBBBBB,
32'h11111111
};
parameter bit [31:0] map_tile14 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000888,
32'h80088CCC,
32'hC88CCCCC,
32'hBCCCCCBC,
32'hBCCCCBBB,
32'hBCCCBBBB,
32'hBBCBBBBB,
32'hBBC9BBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB9BB,
32'hBB3BBBBB,
32'hBBBBBBB9,
32'hBBBBBBBB,
32'hBBBBBBB3,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB33BB9BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB3BBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hB3BBBB3B,
32'h3BBBB9BB,
32'hBBBB3BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h3BBBBB3B,
32'hBBB9BBBB,
32'hBBBBBBBB,
32'h9BBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBB7,
32'hBBBBBBBB,
32'hB9BBB3BB,
32'hBB39BBBB,
32'h3BBBBBBB,
32'hBBBBBBBB,
32'h3BBB9BBB,
32'h7BBBBBBB,
32'hBBB9B9B3,
32'hBB3BBBBB,
32'hBBBBBB3B,
32'hBBBBBB3B,
32'hBBBBBB3B,
32'hB3BBB3BB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBB7B3,
32'hB3B3BBBB,
32'hBBBB3BBB,
32'h579BB7B3,
32'hBBBBBBBB,
32'hB9BBBBBB,
32'hBBBBBBBB,
32'hBB5BBB3B,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h11111111};
parameter bit [31:0] map_tile15 [99:0]='{32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00000000,
32'h00880808,
32'h08CC8C8C,
32'h8CCCCCCB,
32'hCCCCCBBB,
32'hBBCCCBBB,
32'hBBBCBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBB3,
32'hBBB3BBBB,
32'hBBBBBBBB,
32'hB33BB3B3,
32'hBBBBB9BB,
32'h3BBBBBBB,
32'hBBBB9BBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBBB9BBB3,
32'hBB3BBBBB,
32'hB79BBB9B,
32'hBBBB9BBB,
32'hBBBBBB9B,
32'h9B93BBBB,
32'h39BBBBBB,
32'hBBB3BBBB,
32'hBBBBBBBB,
32'hB3BBB3BB,
32'hBBBBBBBB,
32'hBBBBBBB9,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'hBB9BB9BB,
32'hBBBBB3BB,
32'hBBBB9BBB,
32'hBBBB9BBB,
32'h3BBBBBBB,
32'h39BBBBB9,
32'hB9BBBB3B,
32'hBBBBBBBB,
32'hB3BBBBBB,
32'hBBBBBB9B,
32'hBB9BBB9B,
32'hBBBBBBBB,
32'hB5B5BBBB,
32'hBBB597BB,
32'hBB3BBBB7,
32'hBBBBBBB3,
32'hBBBB7BB3,
32'h3BBBBBB9,
32'hBBBBB5BB,
32'hBB3BBBB3,
32'hBBBB9BBB,
32'hBBBBBBB3,
32'h33B7B5BB,
32'hB33BBBB9,
32'hBBBBBBBB,
32'hBBBBBBBB,
32'h11111111
};

logic [511:0]map[99:0];

always_ff @(posedge Clk)
begin
	if(Reset_h)
	begin
map[0]<={map_tile0[0],map_tile1[0],map_tile2[0],map_tile3[0],map_tile4[0],map_tile5[0],map_tile6[0],map_tile7[0],map_tile8[0],map_tile9[0],map_tile10[0],map_tile11[0],map_tile12[0],map_tile13[0],map_tile14[0],map_tile15[0]};
map[1]<={map_tile0[1],map_tile1[1],map_tile2[1],map_tile3[1],map_tile4[1],map_tile5[1],map_tile6[1],map_tile7[1],map_tile8[1],map_tile9[1],map_tile10[1],map_tile11[1],map_tile12[1],map_tile13[1],map_tile14[1],map_tile15[1]};
map[2]<={map_tile0[2],map_tile1[2],map_tile2[2],map_tile3[2],map_tile4[2],map_tile5[2],map_tile6[2],map_tile7[2],map_tile8[2],map_tile9[2],map_tile10[2],map_tile11[2],map_tile12[2],map_tile13[2],map_tile14[2],map_tile15[2]};
map[3]<={map_tile0[3],map_tile1[3],map_tile2[3],map_tile3[3],map_tile4[3],map_tile5[3],map_tile6[3],map_tile7[3],map_tile8[3],map_tile9[3],map_tile10[3],map_tile11[3],map_tile12[3],map_tile13[3],map_tile14[3],map_tile15[3]};
map[4]<={map_tile0[4],map_tile1[4],map_tile2[4],map_tile3[4],map_tile4[4],map_tile5[4],map_tile6[4],map_tile7[4],map_tile8[4],map_tile9[4],map_tile10[4],map_tile11[4],map_tile12[4],map_tile13[4],map_tile14[4],map_tile15[4]};
map[5]<={map_tile0[5],map_tile1[5],map_tile2[5],map_tile3[5],map_tile4[5],map_tile5[5],map_tile6[5],map_tile7[5],map_tile8[5],map_tile9[5],map_tile10[5],map_tile11[5],map_tile12[5],map_tile13[5],map_tile14[5],map_tile15[5]};
map[6]<={map_tile0[6],map_tile1[6],map_tile2[6],map_tile3[6],map_tile4[6],map_tile5[6],map_tile6[6],map_tile7[6],map_tile8[6],map_tile9[6],map_tile10[6],map_tile11[6],map_tile12[6],map_tile13[6],map_tile14[6],map_tile15[6]};
map[7]<={map_tile0[7],map_tile1[7],map_tile2[7],map_tile3[7],map_tile4[7],map_tile5[7],map_tile6[7],map_tile7[7],map_tile8[7],map_tile9[7],map_tile10[7],map_tile11[7],map_tile12[7],map_tile13[7],map_tile14[7],map_tile15[7]};
map[8]<={map_tile0[8],map_tile1[8],map_tile2[8],map_tile3[8],map_tile4[8],map_tile5[8],map_tile6[8],map_tile7[8],map_tile8[8],map_tile9[8],map_tile10[8],map_tile11[8],map_tile12[8],map_tile13[8],map_tile14[8],map_tile15[8]};
map[9]<={map_tile0[9],map_tile1[9],map_tile2[9],map_tile3[9],map_tile4[9],map_tile5[9],map_tile6[9],map_tile7[9],map_tile8[9],map_tile9[9],map_tile10[9],map_tile11[9],map_tile12[9],map_tile13[9],map_tile14[9],map_tile15[9]};
map[10]<={map_tile0[10],map_tile1[10],map_tile2[10],map_tile3[10],map_tile4[10],map_tile5[10],map_tile6[10],map_tile7[10],map_tile8[10],map_tile9[10],map_tile10[10],map_tile11[10],map_tile12[10],map_tile13[10],map_tile14[10],map_tile15[10]};
map[11]<={map_tile0[11],map_tile1[11],map_tile2[11],map_tile3[11],map_tile4[11],map_tile5[11],map_tile6[11],map_tile7[11],map_tile8[11],map_tile9[11],map_tile10[11],map_tile11[11],map_tile12[11],map_tile13[11],map_tile14[11],map_tile15[11]};
map[12]<={map_tile0[12],map_tile1[12],map_tile2[12],map_tile3[12],map_tile4[12],map_tile5[12],map_tile6[12],map_tile7[12],map_tile8[12],map_tile9[12],map_tile10[12],map_tile11[12],map_tile12[12],map_tile13[12],map_tile14[12],map_tile15[12]};
map[13]<={map_tile0[13],map_tile1[13],map_tile2[13],map_tile3[13],map_tile4[13],map_tile5[13],map_tile6[13],map_tile7[13],map_tile8[13],map_tile9[13],map_tile10[13],map_tile11[13],map_tile12[13],map_tile13[13],map_tile14[13],map_tile15[13]};
map[14]<={map_tile0[14],map_tile1[14],map_tile2[14],map_tile3[14],map_tile4[14],map_tile5[14],map_tile6[14],map_tile7[14],map_tile8[14],map_tile9[14],map_tile10[14],map_tile11[14],map_tile12[14],map_tile13[14],map_tile14[14],map_tile15[14]};
map[15]<={map_tile0[15],map_tile1[15],map_tile2[15],map_tile3[15],map_tile4[15],map_tile5[15],map_tile6[15],map_tile7[15],map_tile8[15],map_tile9[15],map_tile10[15],map_tile11[15],map_tile12[15],map_tile13[15],map_tile14[15],map_tile15[15]};
map[16]<={map_tile0[16],map_tile1[16],map_tile2[16],map_tile3[16],map_tile4[16],map_tile5[16],map_tile6[16],map_tile7[16],map_tile8[16],map_tile9[16],map_tile10[16],map_tile11[16],map_tile12[16],map_tile13[16],map_tile14[16],map_tile15[16]};
map[17]<={map_tile0[17],map_tile1[17],map_tile2[17],map_tile3[17],map_tile4[17],map_tile5[17],map_tile6[17],map_tile7[17],map_tile8[17],map_tile9[17],map_tile10[17],map_tile11[17],map_tile12[17],map_tile13[17],map_tile14[17],map_tile15[17]};
map[18]<={map_tile0[18],map_tile1[18],map_tile2[18],map_tile3[18],map_tile4[18],map_tile5[18],map_tile6[18],map_tile7[18],map_tile8[18],map_tile9[18],map_tile10[18],map_tile11[18],map_tile12[18],map_tile13[18],map_tile14[18],map_tile15[18]};
map[19]<={map_tile0[19],map_tile1[19],map_tile2[19],map_tile3[19],map_tile4[19],map_tile5[19],map_tile6[19],map_tile7[19],map_tile8[19],map_tile9[19],map_tile10[19],map_tile11[19],map_tile12[19],map_tile13[19],map_tile14[19],map_tile15[19]};
map[20]<={map_tile0[20],map_tile1[20],map_tile2[20],map_tile3[20],map_tile4[20],map_tile5[20],map_tile6[20],map_tile7[20],map_tile8[20],map_tile9[20],map_tile10[20],map_tile11[20],map_tile12[20],map_tile13[20],map_tile14[20],map_tile15[20]};
map[21]<={map_tile0[21],map_tile1[21],map_tile2[21],map_tile3[21],map_tile4[21],map_tile5[21],map_tile6[21],map_tile7[21],map_tile8[21],map_tile9[21],map_tile10[21],map_tile11[21],map_tile12[21],map_tile13[21],map_tile14[21],map_tile15[21]};
map[22]<={map_tile0[22],map_tile1[22],map_tile2[22],map_tile3[22],map_tile4[22],map_tile5[22],map_tile6[22],map_tile7[22],map_tile8[22],map_tile9[22],map_tile10[22],map_tile11[22],map_tile12[22],map_tile13[22],map_tile14[22],map_tile15[22]};
map[23]<={map_tile0[23],map_tile1[23],map_tile2[23],map_tile3[23],map_tile4[23],map_tile5[23],map_tile6[23],map_tile7[23],map_tile8[23],map_tile9[23],map_tile10[23],map_tile11[23],map_tile12[23],map_tile13[23],map_tile14[23],map_tile15[23]};
map[24]<={map_tile0[24],map_tile1[24],map_tile2[24],map_tile3[24],map_tile4[24],map_tile5[24],map_tile6[24],map_tile7[24],map_tile8[24],map_tile9[24],map_tile10[24],map_tile11[24],map_tile12[24],map_tile13[24],map_tile14[24],map_tile15[24]};
map[25]<={map_tile0[25],map_tile1[25],map_tile2[25],map_tile3[25],map_tile4[25],map_tile5[25],map_tile6[25],map_tile7[25],map_tile8[25],map_tile9[25],map_tile10[25],map_tile11[25],map_tile12[25],map_tile13[25],map_tile14[25],map_tile15[25]};
map[26]<={map_tile0[26],map_tile1[26],map_tile2[26],map_tile3[26],map_tile4[26],map_tile5[26],map_tile6[26],map_tile7[26],map_tile8[26],map_tile9[26],map_tile10[26],map_tile11[26],map_tile12[26],map_tile13[26],map_tile14[26],map_tile15[26]};
map[27]<={map_tile0[27],map_tile1[27],map_tile2[27],map_tile3[27],map_tile4[27],map_tile5[27],map_tile6[27],map_tile7[27],map_tile8[27],map_tile9[27],map_tile10[27],map_tile11[27],map_tile12[27],map_tile13[27],map_tile14[27],map_tile15[27]};
map[28]<={map_tile0[28],map_tile1[28],map_tile2[28],map_tile3[28],map_tile4[28],map_tile5[28],map_tile6[28],map_tile7[28],map_tile8[28],map_tile9[28],map_tile10[28],map_tile11[28],map_tile12[28],map_tile13[28],map_tile14[28],map_tile15[28]};
map[29]<={map_tile0[29],map_tile1[29],map_tile2[29],map_tile3[29],map_tile4[29],map_tile5[29],map_tile6[29],map_tile7[29],map_tile8[29],map_tile9[29],map_tile10[29],map_tile11[29],map_tile12[29],map_tile13[29],map_tile14[29],map_tile15[29]};
map[30]<={map_tile0[30],map_tile1[30],map_tile2[30],map_tile3[30],map_tile4[30],map_tile5[30],map_tile6[30],map_tile7[30],map_tile8[30],map_tile9[30],map_tile10[30],map_tile11[30],map_tile12[30],map_tile13[30],map_tile14[30],map_tile15[30]};
map[31]<={map_tile0[31],map_tile1[31],map_tile2[31],map_tile3[31],map_tile4[31],map_tile5[31],map_tile6[31],map_tile7[31],map_tile8[31],map_tile9[31],map_tile10[31],map_tile11[31],map_tile12[31],map_tile13[31],map_tile14[31],map_tile15[31]};
map[32]<={map_tile0[32],map_tile1[32],map_tile2[32],map_tile3[32],map_tile4[32],map_tile5[32],map_tile6[32],map_tile7[32],map_tile8[32],map_tile9[32],map_tile10[32],map_tile11[32],map_tile12[32],map_tile13[32],map_tile14[32],map_tile15[32]};
map[33]<={map_tile0[33],map_tile1[33],map_tile2[33],map_tile3[33],map_tile4[33],map_tile5[33],map_tile6[33],map_tile7[33],map_tile8[33],map_tile9[33],map_tile10[33],map_tile11[33],map_tile12[33],map_tile13[33],map_tile14[33],map_tile15[33]};
map[34]<={map_tile0[34],map_tile1[34],map_tile2[34],map_tile3[34],map_tile4[34],map_tile5[34],map_tile6[34],map_tile7[34],map_tile8[34],map_tile9[34],map_tile10[34],map_tile11[34],map_tile12[34],map_tile13[34],map_tile14[34],map_tile15[34]};
map[35]<={map_tile0[35],map_tile1[35],map_tile2[35],map_tile3[35],map_tile4[35],map_tile5[35],map_tile6[35],map_tile7[35],map_tile8[35],map_tile9[35],map_tile10[35],map_tile11[35],map_tile12[35],map_tile13[35],map_tile14[35],map_tile15[35]};
map[36]<={map_tile0[36],map_tile1[36],map_tile2[36],map_tile3[36],map_tile4[36],map_tile5[36],map_tile6[36],map_tile7[36],map_tile8[36],map_tile9[36],map_tile10[36],map_tile11[36],map_tile12[36],map_tile13[36],map_tile14[36],map_tile15[36]};
map[37]<={map_tile0[37],map_tile1[37],map_tile2[37],map_tile3[37],map_tile4[37],map_tile5[37],map_tile6[37],map_tile7[37],map_tile8[37],map_tile9[37],map_tile10[37],map_tile11[37],map_tile12[37],map_tile13[37],map_tile14[37],map_tile15[37]};
map[38]<={map_tile0[38],map_tile1[38],map_tile2[38],map_tile3[38],map_tile4[38],map_tile5[38],map_tile6[38],map_tile7[38],map_tile8[38],map_tile9[38],map_tile10[38],map_tile11[38],map_tile12[38],map_tile13[38],map_tile14[38],map_tile15[38]};
map[39]<={map_tile0[39],map_tile1[39],map_tile2[39],map_tile3[39],map_tile4[39],map_tile5[39],map_tile6[39],map_tile7[39],map_tile8[39],map_tile9[39],map_tile10[39],map_tile11[39],map_tile12[39],map_tile13[39],map_tile14[39],map_tile15[39]};
map[40]<={map_tile0[40],map_tile1[40],map_tile2[40],map_tile3[40],map_tile4[40],map_tile5[40],map_tile6[40],map_tile7[40],map_tile8[40],map_tile9[40],map_tile10[40],map_tile11[40],map_tile12[40],map_tile13[40],map_tile14[40],map_tile15[40]};
map[41]<={map_tile0[41],map_tile1[41],map_tile2[41],map_tile3[41],map_tile4[41],map_tile5[41],map_tile6[41],map_tile7[41],map_tile8[41],map_tile9[41],map_tile10[41],map_tile11[41],map_tile12[41],map_tile13[41],map_tile14[41],map_tile15[41]};
map[42]<={map_tile0[42],map_tile1[42],map_tile2[42],map_tile3[42],map_tile4[42],map_tile5[42],map_tile6[42],map_tile7[42],map_tile8[42],map_tile9[42],map_tile10[42],map_tile11[42],map_tile12[42],map_tile13[42],map_tile14[42],map_tile15[42]};
map[43]<={map_tile0[43],map_tile1[43],map_tile2[43],map_tile3[43],map_tile4[43],map_tile5[43],map_tile6[43],map_tile7[43],map_tile8[43],map_tile9[43],map_tile10[43],map_tile11[43],map_tile12[43],map_tile13[43],map_tile14[43],map_tile15[43]};
map[44]<={map_tile0[44],map_tile1[44],map_tile2[44],map_tile3[44],map_tile4[44],map_tile5[44],map_tile6[44],map_tile7[44],map_tile8[44],map_tile9[44],map_tile10[44],map_tile11[44],map_tile12[44],map_tile13[44],map_tile14[44],map_tile15[44]};
map[45]<={map_tile0[45],map_tile1[45],map_tile2[45],map_tile3[45],map_tile4[45],map_tile5[45],map_tile6[45],map_tile7[45],map_tile8[45],map_tile9[45],map_tile10[45],map_tile11[45],map_tile12[45],map_tile13[45],map_tile14[45],map_tile15[45]};
map[46]<={map_tile0[46],map_tile1[46],map_tile2[46],map_tile3[46],map_tile4[46],map_tile5[46],map_tile6[46],map_tile7[46],map_tile8[46],map_tile9[46],map_tile10[46],map_tile11[46],map_tile12[46],map_tile13[46],map_tile14[46],map_tile15[46]};
map[47]<={map_tile0[47],map_tile1[47],map_tile2[47],map_tile3[47],map_tile4[47],map_tile5[47],map_tile6[47],map_tile7[47],map_tile8[47],map_tile9[47],map_tile10[47],map_tile11[47],map_tile12[47],map_tile13[47],map_tile14[47],map_tile15[47]};
map[48]<={map_tile0[48],map_tile1[48],map_tile2[48],map_tile3[48],map_tile4[48],map_tile5[48],map_tile6[48],map_tile7[48],map_tile8[48],map_tile9[48],map_tile10[48],map_tile11[48],map_tile12[48],map_tile13[48],map_tile14[48],map_tile15[48]};
map[49]<={map_tile0[49],map_tile1[49],map_tile2[49],map_tile3[49],map_tile4[49],map_tile5[49],map_tile6[49],map_tile7[49],map_tile8[49],map_tile9[49],map_tile10[49],map_tile11[49],map_tile12[49],map_tile13[49],map_tile14[49],map_tile15[49]};
map[50]<={map_tile0[50],map_tile1[50],map_tile2[50],map_tile3[50],map_tile4[50],map_tile5[50],map_tile6[50],map_tile7[50],map_tile8[50],map_tile9[50],map_tile10[50],map_tile11[50],map_tile12[50],map_tile13[50],map_tile14[50],map_tile15[50]};
map[51]<={map_tile0[51],map_tile1[51],map_tile2[51],map_tile3[51],map_tile4[51],map_tile5[51],map_tile6[51],map_tile7[51],map_tile8[51],map_tile9[51],map_tile10[51],map_tile11[51],map_tile12[51],map_tile13[51],map_tile14[51],map_tile15[51]};
map[52]<={map_tile0[52],map_tile1[52],map_tile2[52],map_tile3[52],map_tile4[52],map_tile5[52],map_tile6[52],map_tile7[52],map_tile8[52],map_tile9[52],map_tile10[52],map_tile11[52],map_tile12[52],map_tile13[52],map_tile14[52],map_tile15[52]};
map[53]<={map_tile0[53],map_tile1[53],map_tile2[53],map_tile3[53],map_tile4[53],map_tile5[53],map_tile6[53],map_tile7[53],map_tile8[53],map_tile9[53],map_tile10[53],map_tile11[53],map_tile12[53],map_tile13[53],map_tile14[53],map_tile15[53]};
map[54]<={map_tile0[54],map_tile1[54],map_tile2[54],map_tile3[54],map_tile4[54],map_tile5[54],map_tile6[54],map_tile7[54],map_tile8[54],map_tile9[54],map_tile10[54],map_tile11[54],map_tile12[54],map_tile13[54],map_tile14[54],map_tile15[54]};
map[55]<={map_tile0[55],map_tile1[55],map_tile2[55],map_tile3[55],map_tile4[55],map_tile5[55],map_tile6[55],map_tile7[55],map_tile8[55],map_tile9[55],map_tile10[55],map_tile11[55],map_tile12[55],map_tile13[55],map_tile14[55],map_tile15[55]};
map[56]<={map_tile0[56],map_tile1[56],map_tile2[56],map_tile3[56],map_tile4[56],map_tile5[56],map_tile6[56],map_tile7[56],map_tile8[56],map_tile9[56],map_tile10[56],map_tile11[56],map_tile12[56],map_tile13[56],map_tile14[56],map_tile15[56]};
map[57]<={map_tile0[57],map_tile1[57],map_tile2[57],map_tile3[57],map_tile4[57],map_tile5[57],map_tile6[57],map_tile7[57],map_tile8[57],map_tile9[57],map_tile10[57],map_tile11[57],map_tile12[57],map_tile13[57],map_tile14[57],map_tile15[57]};
map[58]<={map_tile0[58],map_tile1[58],map_tile2[58],map_tile3[58],map_tile4[58],map_tile5[58],map_tile6[58],map_tile7[58],map_tile8[58],map_tile9[58],map_tile10[58],map_tile11[58],map_tile12[58],map_tile13[58],map_tile14[58],map_tile15[58]};
map[59]<={map_tile0[59],map_tile1[59],map_tile2[59],map_tile3[59],map_tile4[59],map_tile5[59],map_tile6[59],map_tile7[59],map_tile8[59],map_tile9[59],map_tile10[59],map_tile11[59],map_tile12[59],map_tile13[59],map_tile14[59],map_tile15[59]};
map[60]<={map_tile0[60],map_tile1[60],map_tile2[60],map_tile3[60],map_tile4[60],map_tile5[60],map_tile6[60],map_tile7[60],map_tile8[60],map_tile9[60],map_tile10[60],map_tile11[60],map_tile12[60],map_tile13[60],map_tile14[60],map_tile15[60]};
map[61]<={map_tile0[61],map_tile1[61],map_tile2[61],map_tile3[61],map_tile4[61],map_tile5[61],map_tile6[61],map_tile7[61],map_tile8[61],map_tile9[61],map_tile10[61],map_tile11[61],map_tile12[61],map_tile13[61],map_tile14[61],map_tile15[61]};
map[62]<={map_tile0[62],map_tile1[62],map_tile2[62],map_tile3[62],map_tile4[62],map_tile5[62],map_tile6[62],map_tile7[62],map_tile8[62],map_tile9[62],map_tile10[62],map_tile11[62],map_tile12[62],map_tile13[62],map_tile14[62],map_tile15[62]};
map[63]<={map_tile0[63],map_tile1[63],map_tile2[63],map_tile3[63],map_tile4[63],map_tile5[63],map_tile6[63],map_tile7[63],map_tile8[63],map_tile9[63],map_tile10[63],map_tile11[63],map_tile12[63],map_tile13[63],map_tile14[63],map_tile15[63]};
map[64]<={map_tile0[64],map_tile1[64],map_tile2[64],map_tile3[64],map_tile4[64],map_tile5[64],map_tile6[64],map_tile7[64],map_tile8[64],map_tile9[64],map_tile10[64],map_tile11[64],map_tile12[64],map_tile13[64],map_tile14[64],map_tile15[64]};
map[65]<={map_tile0[65],map_tile1[65],map_tile2[65],map_tile3[65],map_tile4[65],map_tile5[65],map_tile6[65],map_tile7[65],map_tile8[65],map_tile9[65],map_tile10[65],map_tile11[65],map_tile12[65],map_tile13[65],map_tile14[65],map_tile15[65]};
map[66]<={map_tile0[66],map_tile1[66],map_tile2[66],map_tile3[66],map_tile4[66],map_tile5[66],map_tile6[66],map_tile7[66],map_tile8[66],map_tile9[66],map_tile10[66],map_tile11[66],map_tile12[66],map_tile13[66],map_tile14[66],map_tile15[66]};
map[67]<={map_tile0[67],map_tile1[67],map_tile2[67],map_tile3[67],map_tile4[67],map_tile5[67],map_tile6[67],map_tile7[67],map_tile8[67],map_tile9[67],map_tile10[67],map_tile11[67],map_tile12[67],map_tile13[67],map_tile14[67],map_tile15[67]};
map[68]<={map_tile0[68],map_tile1[68],map_tile2[68],map_tile3[68],map_tile4[68],map_tile5[68],map_tile6[68],map_tile7[68],map_tile8[68],map_tile9[68],map_tile10[68],map_tile11[68],map_tile12[68],map_tile13[68],map_tile14[68],map_tile15[68]};
map[69]<={map_tile0[69],map_tile1[69],map_tile2[69],map_tile3[69],map_tile4[69],map_tile5[69],map_tile6[69],map_tile7[69],map_tile8[69],map_tile9[69],map_tile10[69],map_tile11[69],map_tile12[69],map_tile13[69],map_tile14[69],map_tile15[69]};
map[70]<={map_tile0[70],map_tile1[70],map_tile2[70],map_tile3[70],map_tile4[70],map_tile5[70],map_tile6[70],map_tile7[70],map_tile8[70],map_tile9[70],map_tile10[70],map_tile11[70],map_tile12[70],map_tile13[70],map_tile14[70],map_tile15[70]};
map[71]<={map_tile0[71],map_tile1[71],map_tile2[71],map_tile3[71],map_tile4[71],map_tile5[71],map_tile6[71],map_tile7[71],map_tile8[71],map_tile9[71],map_tile10[71],map_tile11[71],map_tile12[71],map_tile13[71],map_tile14[71],map_tile15[71]};
map[72]<={map_tile0[72],map_tile1[72],map_tile2[72],map_tile3[72],map_tile4[72],map_tile5[72],map_tile6[72],map_tile7[72],map_tile8[72],map_tile9[72],map_tile10[72],map_tile11[72],map_tile12[72],map_tile13[72],map_tile14[72],map_tile15[72]};
map[73]<={map_tile0[73],map_tile1[73],map_tile2[73],map_tile3[73],map_tile4[73],map_tile5[73],map_tile6[73],map_tile7[73],map_tile8[73],map_tile9[73],map_tile10[73],map_tile11[73],map_tile12[73],map_tile13[73],map_tile14[73],map_tile15[73]};
map[74]<={map_tile0[74],map_tile1[74],map_tile2[74],map_tile3[74],map_tile4[74],map_tile5[74],map_tile6[74],map_tile7[74],map_tile8[74],map_tile9[74],map_tile10[74],map_tile11[74],map_tile12[74],map_tile13[74],map_tile14[74],map_tile15[74]};
map[75]<={map_tile0[75],map_tile1[75],map_tile2[75],map_tile3[75],map_tile4[75],map_tile5[75],map_tile6[75],map_tile7[75],map_tile8[75],map_tile9[75],map_tile10[75],map_tile11[75],map_tile12[75],map_tile13[75],map_tile14[75],map_tile15[75]};
map[76]<={map_tile0[76],map_tile1[76],map_tile2[76],map_tile3[76],map_tile4[76],map_tile5[76],map_tile6[76],map_tile7[76],map_tile8[76],map_tile9[76],map_tile10[76],map_tile11[76],map_tile12[76],map_tile13[76],map_tile14[76],map_tile15[76]};
map[77]<={map_tile0[77],map_tile1[77],map_tile2[77],map_tile3[77],map_tile4[77],map_tile5[77],map_tile6[77],map_tile7[77],map_tile8[77],map_tile9[77],map_tile10[77],map_tile11[77],map_tile12[77],map_tile13[77],map_tile14[77],map_tile15[77]};
map[78]<={map_tile0[78],map_tile1[78],map_tile2[78],map_tile3[78],map_tile4[78],map_tile5[78],map_tile6[78],map_tile7[78],map_tile8[78],map_tile9[78],map_tile10[78],map_tile11[78],map_tile12[78],map_tile13[78],map_tile14[78],map_tile15[78]};
map[79]<={map_tile0[79],map_tile1[79],map_tile2[79],map_tile3[79],map_tile4[79],map_tile5[79],map_tile6[79],map_tile7[79],map_tile8[79],map_tile9[79],map_tile10[79],map_tile11[79],map_tile12[79],map_tile13[79],map_tile14[79],map_tile15[79]};
map[80]<={map_tile0[80],map_tile1[80],map_tile2[80],map_tile3[80],map_tile4[80],map_tile5[80],map_tile6[80],map_tile7[80],map_tile8[80],map_tile9[80],map_tile10[80],map_tile11[80],map_tile12[80],map_tile13[80],map_tile14[80],map_tile15[80]};
map[81]<={map_tile0[81],map_tile1[81],map_tile2[81],map_tile3[81],map_tile4[81],map_tile5[81],map_tile6[81],map_tile7[81],map_tile8[81],map_tile9[81],map_tile10[81],map_tile11[81],map_tile12[81],map_tile13[81],map_tile14[81],map_tile15[81]};
map[82]<={map_tile0[82],map_tile1[82],map_tile2[82],map_tile3[82],map_tile4[82],map_tile5[82],map_tile6[82],map_tile7[82],map_tile8[82],map_tile9[82],map_tile10[82],map_tile11[82],map_tile12[82],map_tile13[82],map_tile14[82],map_tile15[82]};
map[83]<={map_tile0[83],map_tile1[83],map_tile2[83],map_tile3[83],map_tile4[83],map_tile5[83],map_tile6[83],map_tile7[83],map_tile8[83],map_tile9[83],map_tile10[83],map_tile11[83],map_tile12[83],map_tile13[83],map_tile14[83],map_tile15[83]};
map[84]<={map_tile0[84],map_tile1[84],map_tile2[84],map_tile3[84],map_tile4[84],map_tile5[84],map_tile6[84],map_tile7[84],map_tile8[84],map_tile9[84],map_tile10[84],map_tile11[84],map_tile12[84],map_tile13[84],map_tile14[84],map_tile15[84]};
map[85]<={map_tile0[85],map_tile1[85],map_tile2[85],map_tile3[85],map_tile4[85],map_tile5[85],map_tile6[85],map_tile7[85],map_tile8[85],map_tile9[85],map_tile10[85],map_tile11[85],map_tile12[85],map_tile13[85],map_tile14[85],map_tile15[85]};
map[86]<={map_tile0[86],map_tile1[86],map_tile2[86],map_tile3[86],map_tile4[86],map_tile5[86],map_tile6[86],map_tile7[86],map_tile8[86],map_tile9[86],map_tile10[86],map_tile11[86],map_tile12[86],map_tile13[86],map_tile14[86],map_tile15[86]};
map[87]<={map_tile0[87],map_tile1[87],map_tile2[87],map_tile3[87],map_tile4[87],map_tile5[87],map_tile6[87],map_tile7[87],map_tile8[87],map_tile9[87],map_tile10[87],map_tile11[87],map_tile12[87],map_tile13[87],map_tile14[87],map_tile15[87]};
map[88]<={map_tile0[88],map_tile1[88],map_tile2[88],map_tile3[88],map_tile4[88],map_tile5[88],map_tile6[88],map_tile7[88],map_tile8[88],map_tile9[88],map_tile10[88],map_tile11[88],map_tile12[88],map_tile13[88],map_tile14[88],map_tile15[88]};
map[89]<={map_tile0[89],map_tile1[89],map_tile2[89],map_tile3[89],map_tile4[89],map_tile5[89],map_tile6[89],map_tile7[89],map_tile8[89],map_tile9[89],map_tile10[89],map_tile11[89],map_tile12[89],map_tile13[89],map_tile14[89],map_tile15[89]};
map[90]<={map_tile0[90],map_tile1[90],map_tile2[90],map_tile3[90],map_tile4[90],map_tile5[90],map_tile6[90],map_tile7[90],map_tile8[90],map_tile9[90],map_tile10[90],map_tile11[90],map_tile12[90],map_tile13[90],map_tile14[90],map_tile15[90]};
map[91]<={map_tile0[91],map_tile1[91],map_tile2[91],map_tile3[91],map_tile4[91],map_tile5[91],map_tile6[91],map_tile7[91],map_tile8[91],map_tile9[91],map_tile10[91],map_tile11[91],map_tile12[91],map_tile13[91],map_tile14[91],map_tile15[91]};
map[92]<={map_tile0[92],map_tile1[92],map_tile2[92],map_tile3[92],map_tile4[92],map_tile5[92],map_tile6[92],map_tile7[92],map_tile8[92],map_tile9[92],map_tile10[92],map_tile11[92],map_tile12[92],map_tile13[92],map_tile14[92],map_tile15[92]};
map[93]<={map_tile0[93],map_tile1[93],map_tile2[93],map_tile3[93],map_tile4[93],map_tile5[93],map_tile6[93],map_tile7[93],map_tile8[93],map_tile9[93],map_tile10[93],map_tile11[93],map_tile12[93],map_tile13[93],map_tile14[93],map_tile15[93]};
map[94]<={map_tile0[94],map_tile1[94],map_tile2[94],map_tile3[94],map_tile4[94],map_tile5[94],map_tile6[94],map_tile7[94],map_tile8[94],map_tile9[94],map_tile10[94],map_tile11[94],map_tile12[94],map_tile13[94],map_tile14[94],map_tile15[94]};
map[95]<={map_tile0[95],map_tile1[95],map_tile2[95],map_tile3[95],map_tile4[95],map_tile5[95],map_tile6[95],map_tile7[95],map_tile8[95],map_tile9[95],map_tile10[95],map_tile11[95],map_tile12[95],map_tile13[95],map_tile14[95],map_tile15[95]};
map[96]<={map_tile0[96],map_tile1[96],map_tile2[96],map_tile3[96],map_tile4[96],map_tile5[96],map_tile6[96],map_tile7[96],map_tile8[96],map_tile9[96],map_tile10[96],map_tile11[96],map_tile12[96],map_tile13[96],map_tile14[96],map_tile15[96]};
map[97]<={map_tile0[97],map_tile1[97],map_tile2[97],map_tile3[97],map_tile4[97],map_tile5[97],map_tile6[97],map_tile7[97],map_tile8[97],map_tile9[97],map_tile10[97],map_tile11[97],map_tile12[97],map_tile13[97],map_tile14[97],map_tile15[97]};
map[98]<={map_tile0[98],map_tile1[98],map_tile2[98],map_tile3[98],map_tile4[98],map_tile5[98],map_tile6[98],map_tile7[98],map_tile8[98],map_tile9[98],map_tile10[98],map_tile11[98],map_tile12[98],map_tile13[98],map_tile14[98],map_tile15[98]};
map[99]<={map_tile0[99],map_tile1[99],map_tile2[99],map_tile3[99],map_tile4[99],map_tile5[99],map_tile6[99],map_tile7[99],map_tile8[99],map_tile9[99],map_tile10[99],map_tile11[99],map_tile12[99],map_tile13[99],map_tile14[99],map_tile15[99]};
	
	end
	
	else
	begin
	if(operation==2'b01) //dig
	begin
	map[99-changey][4*(128-changex)-1-:4]=4'b0000;
	end
	else if (operation==2'b10) // push
	map[99-changey][4*(128-changex)-1-:4]=push_id;
	end

end

*/

parameter bit [95:0] small_map [99:0]='{
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000000000,
96'h000000000000000000A00000,
96'h00000000000000000AAA0000,
96'h0000000000000000AAEAA000,
96'h088000000000000AAAEAAA00,
96'h8CC888888800000000E00000,
96'hCBCCCCCCCC00088000E00000,
96'hCBCCCBCBCC888CC000E80000,
96'hCBCBBBBBCCCCCCC8888C0008,
96'hBBBBBBBBBBBCCCBCCCCC888C,
96'hBBBBBBBBBBBCBCBBCBBCCCCC,
96'hBBBBBBBBBBBBBBBBCBBBBBCC,
96'h3BBBBBBBBBBBBBBBCBBBBBBB,
96'hBBBBB9BBBBBBBBBBBBBBBBBB,
96'hB3B3B3BBBBBBBBBBBBBBBBBB,
96'hBBBBB7BBBBBBBBB9BBBBBBBB,
96'hBB3BBBBBBBBBB3BBBBBBBBBB,
96'hBBBB9BB3BBBB7BBBB3BBBBB3,
96'hBBBBBBBBB37BBBBBBBBBBBBB,
96'hBBBBBBBBB93BBBBBBB9BB3BB,
96'h73BBBBBBBBBBBBBBBB73BB33,
96'hBBBBB3BBBBB3BBB3B3BBBBBB,
96'hBBBBBBB3BBB9BBBB3BBBBBBB,
96'hBBBBBBBBBBBBBBBBBBBBBBBB,
96'h9BB3BBB7BB7BB9BB9BB7BBBB,
96'hBBBBBB3BBBBBBBB3BBBBBBBB,
96'hBBBBB9BBBBBBBBBBBBBB39BB,
96'hBBBB9BBB7BB3BBB9BBBBBBBB,
96'hB3B3BBBBBBBBBBB3BBBBBBBB,
96'hBBBBBBBB9BB9BBBBBB7BBBBB,
96'hBBBBBBBBBBBBBB9BBBBBBBBB,
96'hBBBBBBBB9BBBB3BBB7BBB7BB,
96'hBBBBBB9BBBBBB3BBBBBBBB3B,
96'hB9BB3B7BB93BB33BBBB9BBB9,
96'hBBBBBBBBBBB5B99BBBBBBBBB,
96'hBBBBBBBBBBBBBB3BBBBBB3BB,
96'hBBBB9BBB3BBBBBBBBBBBBBBB,
96'hBBBBBBB3BBBBBBBBBBBBBBBB,
96'hB5BBBBBBB9BBBBB7BBB75BBB,
96'hBBBB5BBBBBB7BBB3BBB3B3BB,
96'hB9B9BBBB3BB3BBB3BBBBBB7B,
96'hBBBBBBBBBBB3BB99BBBBBBBB,
96'hBB7BBBBBBBBBBBBBBBBB939B,
96'hBBB3BBBB57BBBBBBBBBBBB97,
96'hBBBBBBBBBBBB35BBBBB3BBBB,
96'hB9BBBBBBBB3BBBBBBB3BBBBB,
96'hBBBBBBBBBBBBBBBBBB7BBBBB,
96'hBBBBBBBBBBBBBBBBBBBBBBBB,
96'hBBBBBBBBBBBBBBBBBBBB539B,
96'hB3BBBBBBBB3B7BB3BBBB7BBB,
96'hBB3BBBBB3BB7B7BB3BBBBBBB,
96'h3BBBBBBBB7BBBBBBBBBBBBBB,
96'hB9B5BBBB9BBBBBB79BBBBB3B,
96'h111111111111111111111111

};

logic [95:0] map [99:0];

always_ff @(posedge Clk)
begin
if(Reset_h)
begin
	map[0]<=small_map[0];
map[1]<=small_map[1];
map[2]<=small_map[2];
map[3]<=small_map[3];
map[4]<=small_map[4];
map[5]<=small_map[5];
map[6]<=small_map[6];
map[7]<=small_map[7];
map[8]<=small_map[8];
map[9]<=small_map[9];
map[10]<=small_map[10];
map[11]<=small_map[11];
map[12]<=small_map[12];
map[13]<=small_map[13];
map[14]<=small_map[14];
map[15]<=small_map[15];
map[16]<=small_map[16];
map[17]<=small_map[17];
map[18]<=small_map[18];
map[19]<=small_map[19];
map[20]<=small_map[20];
map[21]<=small_map[21];
map[22]<=small_map[22];
map[23]<=small_map[23];
map[24]<=small_map[24];
map[25]<=small_map[25];
map[26]<=small_map[26];
map[27]<=small_map[27];
map[28]<=small_map[28];
map[29]<=small_map[29];
map[30]<=small_map[30];
map[31]<=small_map[31];
map[32]<=small_map[32];
map[33]<=small_map[33];
map[34]<=small_map[34];
map[35]<=small_map[35];
map[36]<=small_map[36];
map[37]<=small_map[37];
map[38]<=small_map[38];
map[39]<=small_map[39];
map[40]<=small_map[40];
map[41]<=small_map[41];
map[42]<=small_map[42];
map[43]<=small_map[43];
map[44]<=small_map[44];
map[45]<=small_map[45];
map[46]<=small_map[46];
map[47]<=small_map[47];
map[48]<=small_map[48];
map[49]<=small_map[49];
map[50]<=small_map[50];
map[51]<=small_map[51];
map[52]<=small_map[52];
map[53]<=small_map[53];
map[54]<=small_map[54];
map[55]<=small_map[55];
map[56]<=small_map[56];
map[57]<=small_map[57];
map[58]<=small_map[58];
map[59]<=small_map[59];
map[60]<=small_map[60];
map[61]<=small_map[61];
map[62]<=small_map[62];
map[63]<=small_map[63];
map[64]<=small_map[64];
map[65]<=small_map[65];
map[66]<=small_map[66];
map[67]<=small_map[67];
map[68]<=small_map[68];
map[69]<=small_map[69];
map[70]<=small_map[70];
map[71]<=small_map[71];
map[72]<=small_map[72];
map[73]<=small_map[73];
map[74]<=small_map[74];
map[75]<=small_map[75];
map[76]<=small_map[76];
map[77]<=small_map[77];
map[78]<=small_map[78];
map[79]<=small_map[79];
map[80]<=small_map[80];
map[81]<=small_map[81];
map[82]<=small_map[82];
map[83]<=small_map[83];
map[84]<=small_map[84];
map[85]<=small_map[85];
map[86]<=small_map[86];
map[87]<=small_map[87];
map[88]<=small_map[88];
map[89]<=small_map[89];
map[90]<=small_map[90];
map[91]<=small_map[91];
map[92]<=small_map[92];
map[93]<=small_map[93];
map[94]<=small_map[94];
map[95]<=small_map[95];
map[96]<=small_map[96];
map[97]<=small_map[97];
map[98]<=small_map[98];
map[99]<=small_map[99];

end

	else
	begin
	if(operation==2'b01) //dig
	begin
	map[99-changey][4*(24-changex)-1-:4]<=4'b0000;
	end
	else if (operation==2'b10) // push
	map[99-changey][4*(24-changex)-1-:4]<=push_id;
	end

end

assign row_0=map[99-(corner_y+0)][4*(24-corner_x)-1-:64];
assign row_1=map[99-(corner_y+1)][4*(24-corner_x)-1-:64];
assign row_2=map[99-(corner_y+2)][4*(24-corner_x)-1-:64];
assign row_3=map[99-(corner_y+3)][4*(24-corner_x)-1-:64];
assign row_4=map[99-(corner_y+4)][4*(24-corner_x)-1-:64];
assign row_5=map[99-(corner_y+5)][4*(24-corner_x)-1-:64];
assign row_6=map[99-(corner_y+6)][4*(24-corner_x)-1-:64];
assign row_7=map[99-(corner_y+7)][4*(24-corner_x)-1-:64];
assign row_8=map[99-(corner_y+8)][4*(24-corner_x)-1-:64];
assign row_9=map[99-(corner_y+9)][4*(24-corner_x)-1-:64];
assign row_10=map[99-(corner_y+10)][4*(24-corner_x)-1-:64];
assign row_11=map[99-(corner_y+11)][4*(24-corner_x)-1-:64];

endmodule