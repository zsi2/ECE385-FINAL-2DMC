module false_map

(

	input logic [6:0] corner_x,corner_y, // lefttop corner of buffer
	
	output logic [63:0] row_0,row_1,row_2,row_3,row_4,row_5,row_6,row_7,row_8,row_9,row_10,row_11


);

	parameter bit [95:0] false_map [99:0]= '{
	
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000,
96'b000000000000000000000000000000000000000000000000000001000100010001000100010001000100010001000100,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011,
96'b001100110011001100110011001100110011001100110011001100110011001100110011001100110011001100110011	};

assign row_0=false_map[99-(corner_y+0)][4*(24-corner_x)-1-:64];
assign row_1=false_map[99-(corner_y+1)][4*(24-corner_x)-1-:64];
assign row_2=false_map[99-(corner_y+2)][4*(24-corner_x)-1-:64];
assign row_3=false_map[99-(corner_y+3)][4*(24-corner_x)-1-:64];
assign row_4=false_map[99-(corner_y+4)][4*(24-corner_x)-1-:64];
assign row_5=false_map[99-(corner_y+5)][4*(24-corner_x)-1-:64];
assign row_6=false_map[99-(corner_y+6)][4*(24-corner_x)-1-:64];
assign row_7=false_map[99-(corner_y+7)][4*(24-corner_x)-1-:64];
assign row_8=false_map[99-(corner_y+8)][4*(24-corner_x)-1-:64];
assign row_9=false_map[99-(corner_y+9)][4*(24-corner_x)-1-:64];
assign row_10=false_map[99-(corner_y+10)][4*(24-corner_x)-1-:64];
assign row_11=false_map[99-(corner_y+11)][4*(24-corner_x)-1-:64];

endmodule