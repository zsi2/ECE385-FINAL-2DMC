module artrom
(
	input logic [3:0] id,
	
	input logic [5:0] relx,rely,
	
	input logic [6:0] steve_relx,steve_rely,
	
	
	output logic [23:0] rgb,steve_rgb
	

	
);
	parameter bit [23:0] rom_bedrock [1599:0]='{
	
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h000000,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h000000,
24'h000000,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h979797,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757,
24'h575757


		
};

parameter bit [23:0] rom_wood [1599:0]='{

24'h463926,
24'h463926,
24'h695433,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h685332,
24'h685332,
24'h685332,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6d5837,
24'h6d5837,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h463926,
24'h463926,
24'h695433,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h685332,
24'h685332,
24'h685332,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6d5837,
24'h6d5837,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h6f5a39,
24'h6f5a39,
24'h382b18,
24'h382b18,
24'h382b18,
24'h3f321f,
24'h3f321f,
24'h987849,
24'h987849,
24'h987849,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h665130,
24'h99794a,
24'h99794a,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h685332,
24'h685332,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h957546,
24'h957546,
24'h957546,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h6f5a39,
24'h6f5a39,
24'h382b18,
24'h382b18,
24'h382b18,
24'h3f321f,
24'h3f321f,
24'h987849,
24'h987849,
24'h987849,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h665130,
24'h99794a,
24'h99794a,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h685332,
24'h685332,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h957546,
24'h957546,
24'h957546,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h6f5a39,
24'h6f5a39,
24'h382b18,
24'h382b18,
24'h382b18,
24'h3f321f,
24'h3f321f,
24'h987849,
24'h987849,
24'h987849,
24'h413421,
24'h413421,
24'h665130,
24'h665130,
24'h665130,
24'h99794a,
24'h99794a,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h685332,
24'h685332,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h957546,
24'h957546,
24'h957546,
24'h3a2d1a,
24'h3a2d1a,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h644f2e,
24'h644f2e,
24'h413421,
24'h413421,
24'h413421,
24'h685332,
24'h685332,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3e311e,
24'h3e311e,
24'h675231,
24'h675231,
24'h675231,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3a2d1a,
24'h3a2d1a,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h644f2e,
24'h644f2e,
24'h413421,
24'h413421,
24'h413421,
24'h685332,
24'h685332,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3e311e,
24'h3e311e,
24'h675231,
24'h675231,
24'h675231,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h99794a,
24'h99794a,
24'h99794a,
24'h6d5837,
24'h6d5837,
24'h453825,
24'h453825,
24'h453825,
24'h634e2d,
24'h634e2d,
24'h403320,
24'h403320,
24'h403320,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h987849,
24'h3d301d,
24'h3d301d,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h423522,
24'h423522,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6d5837,
24'h6d5837,
24'h453825,
24'h453825,
24'h453825,
24'h634e2d,
24'h634e2d,
24'h403320,
24'h403320,
24'h403320,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h987849,
24'h3d301d,
24'h3d301d,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h423522,
24'h423522,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6d5837,
24'h6d5837,
24'h453825,
24'h453825,
24'h453825,
24'h634e2d,
24'h634e2d,
24'h403320,
24'h403320,
24'h403320,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h987849,
24'h3d301d,
24'h3d301d,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h423522,
24'h423522,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6a5534,
24'h6a5534,
24'h413421,
24'h413421,
24'h413421,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h675231,
24'h6e5938,
24'h6e5938,
24'h423522,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3c2f1c,
24'h3c2f1c,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6a5534,
24'h6a5534,
24'h413421,
24'h413421,
24'h413421,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h675231,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h675231,
24'h6e5938,
24'h6e5938,
24'h423522,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3c2f1c,
24'h3c2f1c,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h6c5736,
24'h6c5736,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h665130,
24'h665130,
24'h665130,
24'h9a7a4b,
24'h9a7a4b,
24'h685332,
24'h685332,
24'h685332,
24'h665130,
24'h665130,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6b5635,
24'h6b5635,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h695433,
24'h695433,
24'h8f6f40,
24'h8f6f40,
24'h8f6f40,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h675231,
24'h675231,
24'h675231,
24'h6c5736,
24'h6c5736,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h665130,
24'h665130,
24'h665130,
24'h9a7a4b,
24'h9a7a4b,
24'h685332,
24'h685332,
24'h685332,
24'h665130,
24'h665130,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6b5635,
24'h6b5635,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h695433,
24'h695433,
24'h8f6f40,
24'h8f6f40,
24'h8f6f40,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h675231,
24'h675231,
24'h675231,
24'h6c5736,
24'h6c5736,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h665130,
24'h665130,
24'h665130,
24'h9a7a4b,
24'h9a7a4b,
24'h685332,
24'h685332,
24'h685332,
24'h665130,
24'h665130,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6b5635,
24'h6b5635,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h695433,
24'h695433,
24'h8f6f40,
24'h8f6f40,
24'h8f6f40,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h675231,
24'h675231,
24'h675231,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h624d2c,
24'h624d2c,
24'h624d2c,
24'h685332,
24'h685332,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h917142,
24'h917142,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h7c623e,
24'h7c623e,
24'h59472c,
24'h59472c,
24'h59472c,
24'h372a17,
24'h372a17,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h624d2c,
24'h624d2c,
24'h624d2c,
24'h685332,
24'h685332,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h917142,
24'h917142,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h7c623e,
24'h7c623e,
24'h59472c,
24'h59472c,
24'h59472c,
24'h372a17,
24'h372a17,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3e311e,
24'h3e311e,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h413421,
24'h413421,
24'h413421,
24'h99794a,
24'h99794a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h4c3d26,
24'h665130,
24'h665130,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3e311e,
24'h3e311e,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h413421,
24'h413421,
24'h413421,
24'h99794a,
24'h99794a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h4c3d26,
24'h665130,
24'h665130,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h3e311e,
24'h3e311e,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h9b7b4c,
24'h9b7b4c,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h9a7a4b,
24'h9a7a4b,
24'h413421,
24'h413421,
24'h413421,
24'h99794a,
24'h99794a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h4c3d26,
24'h665130,
24'h665130,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h695433,
24'h695433,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3f321f,
24'h3f321f,
24'h705b3a,
24'h705b3a,
24'h705b3a,
24'h947445,
24'h947445,
24'h413421,
24'h413421,
24'h413421,
24'h695433,
24'h695433,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h423522,
24'h423522,
24'h423522,
24'h937344,
24'h937344,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h6c5736,
24'h6c5736,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h3f321f,
24'h3f321f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h99794a,
24'h99794a,
24'h99794a,
24'h3f321f,
24'h3f321f,
24'h705b3a,
24'h705b3a,
24'h705b3a,
24'h947445,
24'h947445,
24'h413421,
24'h413421,
24'h413421,
24'h695433,
24'h695433,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h423522,
24'h423522,
24'h423522,
24'h937344,
24'h937344,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h6c5736,
24'h6c5736,
24'h6b5635,
24'h6b5635,
24'h6b5635,
24'h3f321f,
24'h3f321f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h463926,
24'h463926,
24'h675231,
24'h675231,
24'h675231,
24'h6d5837,
24'h6d5837,
24'h947445,
24'h947445,
24'h947445,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h392c19,
24'h392c19,
24'h392c19,
24'h957546,
24'h957546,
24'h423522,
24'h423522,
24'h423522,
24'h6b5635,
24'h6b5635,
24'h957546,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h463926,
24'h463926,
24'h675231,
24'h675231,
24'h675231,
24'h6d5837,
24'h6d5837,
24'h947445,
24'h947445,
24'h947445,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h392c19,
24'h392c19,
24'h392c19,
24'h957546,
24'h957546,
24'h423522,
24'h423522,
24'h423522,
24'h6b5635,
24'h6b5635,
24'h957546,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h695433,
24'h695433,
24'h9c7c4d,
24'h9c7c4d,
24'h9c7c4d,
24'h463926,
24'h463926,
24'h675231,
24'h675231,
24'h675231,
24'h6d5837,
24'h6d5837,
24'h947445,
24'h947445,
24'h947445,
24'h423522,
24'h423522,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h392c19,
24'h392c19,
24'h392c19,
24'h957546,
24'h957546,
24'h423522,
24'h423522,
24'h423522,
24'h6b5635,
24'h6b5635,
24'h957546,
24'h957546,
24'h957546,
24'h413421,
24'h413421,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h453825,
24'h453825,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h675231,
24'h675231,
24'h967647,
24'h967647,
24'h967647,
24'h3a2d1a,
24'h3a2d1a,
24'h644f2e,
24'h644f2e,
24'h644f2e,
24'h3e311e,
24'h3e311e,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9f7f50,
24'h9f7f50,
24'h403320,
24'h403320,
24'h403320,
24'h6a5534,
24'h6a5534,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h433623,
24'h433623,
24'h957546,
24'h957546,
24'h957546,
24'h453825,
24'h453825,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h403320,
24'h403320,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h675231,
24'h675231,
24'h967647,
24'h967647,
24'h967647,
24'h3a2d1a,
24'h3a2d1a,
24'h644f2e,
24'h644f2e,
24'h644f2e,
24'h3e311e,
24'h3e311e,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9f7f50,
24'h9f7f50,
24'h403320,
24'h403320,
24'h403320,
24'h6a5534,
24'h6a5534,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h433623,
24'h433623,
24'h957546,
24'h957546,
24'h957546,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h675231,
24'h675231,
24'h675231,
24'h6f5a39,
24'h6f5a39,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h423522,
24'h423522,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9d7d4e,
24'h9d7d4e,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h675231,
24'h675231,
24'h675231,
24'h6f5a39,
24'h6f5a39,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h423522,
24'h423522,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9d7d4e,
24'h9d7d4e,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3e311e,
24'h3e311e,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3f321f,
24'h3f321f,
24'h675231,
24'h675231,
24'h675231,
24'h6f5a39,
24'h6f5a39,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h423522,
24'h423522,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h5e4b2f,
24'h5e4b2f,
24'h5e4b2f,
24'h9d7d4e,
24'h9d7d4e,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6c5736,
24'h6c5736,
24'h977748,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h9b7b4c,
24'h9b7b4c,
24'h9b7b4c,
24'h3b2e1b,
24'h3b2e1b,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h392c19,
24'h392c19,
24'h665130,
24'h665130,
24'h665130,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h6a5534,
24'h6a5534,
24'h624d2c,
24'h624d2c,
24'h624d2c,
24'h403320,
24'h403320,
24'h987849,
24'h987849,
24'h987849,
24'h3b2e1b,
24'h3b2e1b,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h392c19,
24'h392c19,
24'h665130,
24'h665130,
24'h665130,
24'h6b5635,
24'h6b5635,
24'h9a7a4b,
24'h9a7a4b,
24'h9a7a4b,
24'h382b18,
24'h382b18,
24'h6a5534,
24'h6a5534,
24'h6a5534,
24'h3f321f,
24'h3f321f,
24'h65502f,
24'h65502f,
24'h65502f,
24'h977748,
24'h977748,
24'h3c2f1c,
24'h3c2f1c,
24'h3c2f1c,
24'h6a5534,
24'h6a5534,
24'h624d2c,
24'h624d2c,
24'h624d2c,
24'h403320,
24'h403320,
24'h987849,
24'h987849,
24'h987849,
24'h413421,
24'h413421,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6d5837,
24'h6d5837,
24'h634e2d,
24'h634e2d,
24'h634e2d,
24'h675231,
24'h675231,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6a5534,
24'h6a5534,
24'h947445,
24'h947445,
24'h947445,
24'h9c7c4d,
24'h9c7c4d,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h413421,
24'h413421,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6d5837,
24'h6d5837,
24'h634e2d,
24'h634e2d,
24'h634e2d,
24'h675231,
24'h675231,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6a5534,
24'h6a5534,
24'h947445,
24'h947445,
24'h947445,
24'h9c7c4d,
24'h9c7c4d,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h413421,
24'h413421,
24'h6d5837,
24'h6d5837,
24'h6d5837,
24'h5e4b2f,
24'h5e4b2f,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h6e5938,
24'h6e5938,
24'h6e5938,
24'h6d5837,
24'h6d5837,
24'h634e2d,
24'h634e2d,
24'h634e2d,
24'h675231,
24'h675231,
24'h3d301d,
24'h3d301d,
24'h3d301d,
24'h6a5534,
24'h6a5534,
24'h947445,
24'h947445,
24'h947445,
24'h9c7c4d,
24'h9c7c4d,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h3a2d1a,
24'h675231,
24'h675231,
24'h675231,
24'h977748,
24'h977748,
24'h403320,
24'h403320,
24'h403320,
24'h6b5635,
24'h6b5635,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h927243,
24'h927243,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3b2e1b,
24'h3b2e1b,
24'h3b2e1b,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3d301d,
24'h3d301d,
24'h675231,
24'h675231,
24'h675231,
24'h3a2d1a,
24'h3a2d1a,
24'h675231,
24'h675231,
24'h675231,
24'h977748,
24'h977748,
24'h403320,
24'h403320,
24'h403320,
24'h6b5635,
24'h6b5635,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h4c3d26,
24'h4c3d26,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h927243,
24'h927243,
24'h685332,
24'h685332,
24'h685332,
24'h987849,
24'h987849,
24'h3b2e1b,
24'h3b2e1b,
24'h3b2e1b,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h3d301d,
24'h3d301d,
24'h675231,
24'h675231,
24'h675231,
24'h5e4b2f,
24'h5e4b2f,
24'h685332,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h644f2e,
24'h644f2e,
24'h695433,
24'h695433,
24'h695433,
24'h685332,
24'h685332,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h372a17,
24'h372a17,
24'h372a17,
24'h675231,
24'h675231,
24'h695433,
24'h695433,
24'h695433,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h5e4b2f,
24'h5e4b2f,
24'h685332,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h644f2e,
24'h644f2e,
24'h695433,
24'h695433,
24'h695433,
24'h685332,
24'h685332,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h372a17,
24'h372a17,
24'h372a17,
24'h675231,
24'h675231,
24'h695433,
24'h695433,
24'h695433,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e,
24'h5e4b2f,
24'h5e4b2f,
24'h685332,
24'h685332,
24'h685332,
24'h7c623e,
24'h7c623e,
24'h3e311e,
24'h3e311e,
24'h3e311e,
24'h644f2e,
24'h644f2e,
24'h695433,
24'h695433,
24'h695433,
24'h685332,
24'h685332,
24'h403320,
24'h403320,
24'h403320,
24'h695433,
24'h695433,
24'h6c5736,
24'h6c5736,
24'h6c5736,
24'h675231,
24'h675231,
24'h372a17,
24'h372a17,
24'h372a17,
24'h675231,
24'h675231,
24'h695433,
24'h695433,
24'h695433,
24'h65502f,
24'h65502f,
24'h7c623e,
24'h7c623e,
24'h7c623e




};

parameter bit [23:0] rom_stone [1599:0]='{

24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h808080,
24'h808080,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h808080,
24'h808080,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h808080,
24'h808080,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h686868,
24'h686868,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h686868,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h686868,
24'h686868,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h8f8f8f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h747474,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f,
24'h7f7f7f





};

parameter bit [23:0] rom_dirt [1599:0]='{


24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h979797,
24'h979797,
24'h979797,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h979797,
24'h979797,
24'h979797,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'hb9855c,
24'h79553a,
24'h79553a,
24'h79553a,
24'h79553a




};

parameter bit [23:0] rom_steve [3199:0] ='{

24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h1b1004,
24'h1b1004,
24'h1b1004,
24'h170d01,
24'h170d01,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h100800,
24'h100800,
24'h0d0600,
24'h0d0600,
24'h0d0600,
24'h100800,
24'h100800,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h1b1004,
24'h1b1004,
24'h1b1004,
24'h170d01,
24'h170d01,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h100800,
24'h100800,
24'h0d0600,
24'h0d0600,
24'h0d0600,
24'h100800,
24'h100800,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h1b1004,
24'h1b1004,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h1b1004,
24'h1b1004,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h170d01,
24'h1b1004,
24'h1b1004,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h271a0c,
24'h1a1003,
24'h1a1003,
24'h1a1003,
24'h170d01,
24'h170d01,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h956f5a,
24'h956f5a,
24'h936551,
24'h936551,
24'h936551,
24'h946b57,
24'h946b57,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h211508,
24'h211508,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h956f5a,
24'h956f5a,
24'h936551,
24'h936551,
24'h936551,
24'h946b57,
24'h946b57,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h211508,
24'h211508,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h170d01,
24'h170d01,
24'h170d01,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h956f5a,
24'h956f5a,
24'h936551,
24'h936551,
24'h936551,
24'h946b57,
24'h946b57,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h211508,
24'h211508,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h915c48,
24'h915c48,
24'h915c48,
24'h946752,
24'h946752,
24'h915c48,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h936551,
24'h936551,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h915c48,
24'h915c48,
24'h915c48,
24'h946752,
24'h946752,
24'h915c48,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h8f5944,
24'h8f5944,
24'h8f5944,
24'h936551,
24'h936551,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'h8c543f,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h946752,
24'h946752,
24'h946752,
24'hffffff,
24'hffffff,
24'h312877,
24'h312877,
24'h312877,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h312877,
24'h312877,
24'hffffff,
24'hffffff,
24'hffffff,
24'h915c48,
24'h915c48,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h946752,
24'h946752,
24'h946752,
24'hffffff,
24'hffffff,
24'h312877,
24'h312877,
24'h312877,
24'h915c48,
24'h915c48,
24'h936551,
24'h936551,
24'h936551,
24'h312877,
24'h312877,
24'hffffff,
24'hffffff,
24'hffffff,
24'h915c48,
24'h915c48,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h7b4435,
24'h7b4435,
24'h7b4435,
24'h8b5441,
24'h8b5441,
24'h936551,
24'h936551,
24'h936551,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h936551,
24'h936551,
24'h8d5441,
24'h8d5441,
24'h8d5441,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h7b4435,
24'h7b4435,
24'h7b4435,
24'h8b5441,
24'h8b5441,
24'h936551,
24'h936551,
24'h936551,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h936551,
24'h936551,
24'h8d5441,
24'h8d5441,
24'h8d5441,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h7b4435,
24'h7b4435,
24'h7b4435,
24'h8b5441,
24'h8b5441,
24'h936551,
24'h936551,
24'h936551,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h6b3b2e,
24'h936551,
24'h936551,
24'h8d5441,
24'h8d5441,
24'h8d5441,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h7b4435,
24'h7b4435,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h713b2d,
24'h713b2d,
24'h713b2d,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h7b4435,
24'h7b4435,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h713b2d,
24'h713b2d,
24'h713b2d,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h7b4435,
24'h7b4435,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h61362c,
24'h713b2d,
24'h713b2d,
24'h713b2d,
24'h65372c,
24'h65372c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h764031,
24'h764031,
24'h764031,
24'h764031,
24'h764031,
24'h6a3a2d,
24'h6a3a2d,
24'h6a3a2d,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h60362c,
24'h60362c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h6a372b,
24'h764031,
24'h764031,
24'h764031,
24'h764031,
24'h764031,
24'h6a3a2d,
24'h6a3a2d,
24'h6a3a2d,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h733d2f,
24'h60362c,
24'h60362c,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h905944,
24'h905944,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h905944,
24'h905944,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h008282,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h854837,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h008282,
24'h008282,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h007e7e,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h008b8b,
24'h008b8b,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h009090,
24'h009090,
24'h009090,
24'h007e7e,
24'h007e7e,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h007e7e,
24'h007e7e,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h905944,
24'h936551,
24'h936551,
24'h936551,
24'h905944,
24'h905944,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h312877,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'h3a3088,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'h585858,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff,
24'hffffff



};

	
always_comb
begin
 if(rely<40&relx<40)	
 begin
	if(id==4'b0001)
		rgb= rom_bedrock[rely*40+relx];
	else if(id==4'b0010)
		rgb= rom_wood [rely*40+relx];
	else if(id==4'b0011)
		rgb= rom_stone [rely*40+relx];
	else if(id==4'b0100)
		rgb= rom_dirt [rely*40+relx];
	else
		rgb=24'b0;
 end
 else
 
 rgb=24'b0;
 
end

always_comb
begin
	if((steve_relx!=6'b0)&(steve_rely!=6'b0))
	begin
		steve_rgb=rom_steve[(79-steve_rely)*40+steve_relx];
	end
	
	else
		steve_rgb=24'hd2e6ff;
end







endmodule